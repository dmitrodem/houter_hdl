library ieee;
use ieee.std_logic_1164.all;

entity SpaceWireRouterIPCRCRom is
  port (
    clock   : in  std_logic;
    address : in  std_logic_vector (8 downto 0);
    readData    : out std_logic_vector (7 downto 0));
end entity SpaceWireRouterIPCRCRom;

architecture rtl of SpaceWireRouterIPCRCRom is

  signal romdata : std_logic_vector (readData'range);

begin  -- architecture rtl

  comb : process (address) is
  begin  -- process comb
    case address is
      when "000000000" => romdata <= x"00";
      when "000000001" => romdata <= x"07";
      when "000000010" => romdata <= x"0e";
      when "000000011" => romdata <= x"09";
      when "000000100" => romdata <= x"1c";
      when "000000101" => romdata <= x"1b";
      when "000000110" => romdata <= x"12";
      when "000000111" => romdata <= x"15";
      when "000001000" => romdata <= x"38";
      when "000001001" => romdata <= x"3f";
      when "000001010" => romdata <= x"36";
      when "000001011" => romdata <= x"31";
      when "000001100" => romdata <= x"24";
      when "000001101" => romdata <= x"23";
      when "000001110" => romdata <= x"2a";
      when "000001111" => romdata <= x"2d";
      when "000010000" => romdata <= x"70";
      when "000010001" => romdata <= x"77";
      when "000010010" => romdata <= x"7e";
      when "000010011" => romdata <= x"79";
      when "000010100" => romdata <= x"6c";
      when "000010101" => romdata <= x"6b";
      when "000010110" => romdata <= x"62";
      when "000010111" => romdata <= x"65";
      when "000011000" => romdata <= x"48";
      when "000011001" => romdata <= x"4f";
      when "000011010" => romdata <= x"46";
      when "000011011" => romdata <= x"41";
      when "000011100" => romdata <= x"54";
      when "000011101" => romdata <= x"53";
      when "000011110" => romdata <= x"5a";
      when "000011111" => romdata <= x"5d";
      when "000100000" => romdata <= x"e0";
      when "000100001" => romdata <= x"e7";
      when "000100010" => romdata <= x"ee";
      when "000100011" => romdata <= x"e9";
      when "000100100" => romdata <= x"fc";
      when "000100101" => romdata <= x"fb";
      when "000100110" => romdata <= x"f2";
      when "000100111" => romdata <= x"f5";
      when "000101000" => romdata <= x"d8";
      when "000101001" => romdata <= x"df";
      when "000101010" => romdata <= x"d6";
      when "000101011" => romdata <= x"d1";
      when "000101100" => romdata <= x"c4";
      when "000101101" => romdata <= x"c3";
      when "000101110" => romdata <= x"ca";
      when "000101111" => romdata <= x"cd";
      when "000110000" => romdata <= x"90";
      when "000110001" => romdata <= x"97";
      when "000110010" => romdata <= x"9e";
      when "000110011" => romdata <= x"99";
      when "000110100" => romdata <= x"8c";
      when "000110101" => romdata <= x"8b";
      when "000110110" => romdata <= x"82";
      when "000110111" => romdata <= x"85";
      when "000111000" => romdata <= x"a8";
      when "000111001" => romdata <= x"af";
      when "000111010" => romdata <= x"a6";
      when "000111011" => romdata <= x"a1";
      when "000111100" => romdata <= x"b4";
      when "000111101" => romdata <= x"b3";
      when "000111110" => romdata <= x"ba";
      when "000111111" => romdata <= x"bd";
      when "001000000" => romdata <= x"c7";
      when "001000001" => romdata <= x"c0";
      when "001000010" => romdata <= x"c9";
      when "001000011" => romdata <= x"ce";
      when "001000100" => romdata <= x"db";
      when "001000101" => romdata <= x"dc";
      when "001000110" => romdata <= x"d5";
      when "001000111" => romdata <= x"d2";
      when "001001000" => romdata <= x"ff";
      when "001001001" => romdata <= x"f8";
      when "001001010" => romdata <= x"f1";
      when "001001011" => romdata <= x"f6";
      when "001001100" => romdata <= x"e3";
      when "001001101" => romdata <= x"e4";
      when "001001110" => romdata <= x"ed";
      when "001001111" => romdata <= x"ea";
      when "001010000" => romdata <= x"b7";
      when "001010001" => romdata <= x"b0";
      when "001010010" => romdata <= x"b9";
      when "001010011" => romdata <= x"be";
      when "001010100" => romdata <= x"ab";
      when "001010101" => romdata <= x"ac";
      when "001010110" => romdata <= x"a5";
      when "001010111" => romdata <= x"a2";
      when "001011000" => romdata <= x"8f";
      when "001011001" => romdata <= x"88";
      when "001011010" => romdata <= x"81";
      when "001011011" => romdata <= x"86";
      when "001011100" => romdata <= x"93";
      when "001011101" => romdata <= x"94";
      when "001011110" => romdata <= x"9d";
      when "001011111" => romdata <= x"9a";
      when "001100000" => romdata <= x"27";
      when "001100001" => romdata <= x"20";
      when "001100010" => romdata <= x"29";
      when "001100011" => romdata <= x"2e";
      when "001100100" => romdata <= x"3b";
      when "001100101" => romdata <= x"3c";
      when "001100110" => romdata <= x"35";
      when "001100111" => romdata <= x"32";
      when "001101000" => romdata <= x"1f";
      when "001101001" => romdata <= x"18";
      when "001101010" => romdata <= x"11";
      when "001101011" => romdata <= x"16";
      when "001101100" => romdata <= x"03";
      when "001101101" => romdata <= x"04";
      when "001101110" => romdata <= x"0d";
      when "001101111" => romdata <= x"0a";
      when "001110000" => romdata <= x"57";
      when "001110001" => romdata <= x"50";
      when "001110010" => romdata <= x"59";
      when "001110011" => romdata <= x"5e";
      when "001110100" => romdata <= x"4b";
      when "001110101" => romdata <= x"4c";
      when "001110110" => romdata <= x"45";
      when "001110111" => romdata <= x"42";
      when "001111000" => romdata <= x"6f";
      when "001111001" => romdata <= x"68";
      when "001111010" => romdata <= x"61";
      when "001111011" => romdata <= x"66";
      when "001111100" => romdata <= x"73";
      when "001111101" => romdata <= x"74";
      when "001111110" => romdata <= x"7d";
      when "001111111" => romdata <= x"7a";
      when "010000000" => romdata <= x"89";
      when "010000001" => romdata <= x"8e";
      when "010000010" => romdata <= x"87";
      when "010000011" => romdata <= x"80";
      when "010000100" => romdata <= x"95";
      when "010000101" => romdata <= x"92";
      when "010000110" => romdata <= x"9b";
      when "010000111" => romdata <= x"9c";
      when "010001000" => romdata <= x"b1";
      when "010001001" => romdata <= x"b6";
      when "010001010" => romdata <= x"bf";
      when "010001011" => romdata <= x"b8";
      when "010001100" => romdata <= x"ad";
      when "010001101" => romdata <= x"aa";
      when "010001110" => romdata <= x"a3";
      when "010001111" => romdata <= x"a4";
      when "010010000" => romdata <= x"f9";
      when "010010001" => romdata <= x"fe";
      when "010010010" => romdata <= x"f7";
      when "010010011" => romdata <= x"f0";
      when "010010100" => romdata <= x"e5";
      when "010010101" => romdata <= x"e2";
      when "010010110" => romdata <= x"eb";
      when "010010111" => romdata <= x"ec";
      when "010011000" => romdata <= x"c1";
      when "010011001" => romdata <= x"c6";
      when "010011010" => romdata <= x"cf";
      when "010011011" => romdata <= x"c8";
      when "010011100" => romdata <= x"dd";
      when "010011101" => romdata <= x"da";
      when "010011110" => romdata <= x"d3";
      when "010011111" => romdata <= x"d4";
      when "010100000" => romdata <= x"69";
      when "010100001" => romdata <= x"6e";
      when "010100010" => romdata <= x"67";
      when "010100011" => romdata <= x"60";
      when "010100100" => romdata <= x"75";
      when "010100101" => romdata <= x"72";
      when "010100110" => romdata <= x"7b";
      when "010100111" => romdata <= x"7c";
      when "010101000" => romdata <= x"51";
      when "010101001" => romdata <= x"56";
      when "010101010" => romdata <= x"5f";
      when "010101011" => romdata <= x"58";
      when "010101100" => romdata <= x"4d";
      when "010101101" => romdata <= x"4a";
      when "010101110" => romdata <= x"43";
      when "010101111" => romdata <= x"44";
      when "010110000" => romdata <= x"19";
      when "010110001" => romdata <= x"1e";
      when "010110010" => romdata <= x"17";
      when "010110011" => romdata <= x"10";
      when "010110100" => romdata <= x"05";
      when "010110101" => romdata <= x"02";
      when "010110110" => romdata <= x"0b";
      when "010110111" => romdata <= x"0c";
      when "010111000" => romdata <= x"21";
      when "010111001" => romdata <= x"26";
      when "010111010" => romdata <= x"2f";
      when "010111011" => romdata <= x"28";
      when "010111100" => romdata <= x"3d";
      when "010111101" => romdata <= x"3a";
      when "010111110" => romdata <= x"33";
      when "010111111" => romdata <= x"34";
      when "011000000" => romdata <= x"4e";
      when "011000001" => romdata <= x"49";
      when "011000010" => romdata <= x"40";
      when "011000011" => romdata <= x"47";
      when "011000100" => romdata <= x"52";
      when "011000101" => romdata <= x"55";
      when "011000110" => romdata <= x"5c";
      when "011000111" => romdata <= x"5b";
      when "011001000" => romdata <= x"76";
      when "011001001" => romdata <= x"71";
      when "011001010" => romdata <= x"78";
      when "011001011" => romdata <= x"7f";
      when "011001100" => romdata <= x"6a";
      when "011001101" => romdata <= x"6d";
      when "011001110" => romdata <= x"64";
      when "011001111" => romdata <= x"63";
      when "011010000" => romdata <= x"3e";
      when "011010001" => romdata <= x"39";
      when "011010010" => romdata <= x"30";
      when "011010011" => romdata <= x"37";
      when "011010100" => romdata <= x"22";
      when "011010101" => romdata <= x"25";
      when "011010110" => romdata <= x"2c";
      when "011010111" => romdata <= x"2b";
      when "011011000" => romdata <= x"06";
      when "011011001" => romdata <= x"01";
      when "011011010" => romdata <= x"08";
      when "011011011" => romdata <= x"0f";
      when "011011100" => romdata <= x"1a";
      when "011011101" => romdata <= x"1d";
      when "011011110" => romdata <= x"14";
      when "011011111" => romdata <= x"13";
      when "011100000" => romdata <= x"ae";
      when "011100001" => romdata <= x"a9";
      when "011100010" => romdata <= x"a0";
      when "011100011" => romdata <= x"a7";
      when "011100100" => romdata <= x"b2";
      when "011100101" => romdata <= x"b5";
      when "011100110" => romdata <= x"bc";
      when "011100111" => romdata <= x"bb";
      when "011101000" => romdata <= x"96";
      when "011101001" => romdata <= x"91";
      when "011101010" => romdata <= x"98";
      when "011101011" => romdata <= x"9f";
      when "011101100" => romdata <= x"8a";
      when "011101101" => romdata <= x"8d";
      when "011101110" => romdata <= x"84";
      when "011101111" => romdata <= x"83";
      when "011110000" => romdata <= x"de";
      when "011110001" => romdata <= x"d9";
      when "011110010" => romdata <= x"d0";
      when "011110011" => romdata <= x"d7";
      when "011110100" => romdata <= x"c2";
      when "011110101" => romdata <= x"c5";
      when "011110110" => romdata <= x"cc";
      when "011110111" => romdata <= x"cb";
      when "011111000" => romdata <= x"e6";
      when "011111001" => romdata <= x"e1";
      when "011111010" => romdata <= x"e8";
      when "011111011" => romdata <= x"ef";
      when "011111100" => romdata <= x"fa";
      when "011111101" => romdata <= x"fd";
      when "011111110" => romdata <= x"f4";
      when "011111111" => romdata <= x"f3";
      when "100000000" => romdata <= x"00";
      when "100000001" => romdata <= x"91";
      when "100000010" => romdata <= x"e3";
      when "100000011" => romdata <= x"72";
      when "100000100" => romdata <= x"07";
      when "100000101" => romdata <= x"96";
      when "100000110" => romdata <= x"e4";
      when "100000111" => romdata <= x"75";
      when "100001000" => romdata <= x"0e";
      when "100001001" => romdata <= x"9f";
      when "100001010" => romdata <= x"ed";
      when "100001011" => romdata <= x"7c";
      when "100001100" => romdata <= x"09";
      when "100001101" => romdata <= x"98";
      when "100001110" => romdata <= x"ea";
      when "100001111" => romdata <= x"7b";
      when "100010000" => romdata <= x"1c";
      when "100010001" => romdata <= x"8d";
      when "100010010" => romdata <= x"ff";
      when "100010011" => romdata <= x"6e";
      when "100010100" => romdata <= x"1b";
      when "100010101" => romdata <= x"8a";
      when "100010110" => romdata <= x"f8";
      when "100010111" => romdata <= x"69";
      when "100011000" => romdata <= x"12";
      when "100011001" => romdata <= x"83";
      when "100011010" => romdata <= x"f1";
      when "100011011" => romdata <= x"60";
      when "100011100" => romdata <= x"15";
      when "100011101" => romdata <= x"84";
      when "100011110" => romdata <= x"f6";
      when "100011111" => romdata <= x"67";
      when "100100000" => romdata <= x"38";
      when "100100001" => romdata <= x"a9";
      when "100100010" => romdata <= x"db";
      when "100100011" => romdata <= x"4a";
      when "100100100" => romdata <= x"3f";
      when "100100101" => romdata <= x"ae";
      when "100100110" => romdata <= x"dc";
      when "100100111" => romdata <= x"4d";
      when "100101000" => romdata <= x"36";
      when "100101001" => romdata <= x"a7";
      when "100101010" => romdata <= x"d5";
      when "100101011" => romdata <= x"44";
      when "100101100" => romdata <= x"31";
      when "100101101" => romdata <= x"a0";
      when "100101110" => romdata <= x"d2";
      when "100101111" => romdata <= x"43";
      when "100110000" => romdata <= x"24";
      when "100110001" => romdata <= x"b5";
      when "100110010" => romdata <= x"c7";
      when "100110011" => romdata <= x"56";
      when "100110100" => romdata <= x"23";
      when "100110101" => romdata <= x"b2";
      when "100110110" => romdata <= x"c0";
      when "100110111" => romdata <= x"51";
      when "100111000" => romdata <= x"2a";
      when "100111001" => romdata <= x"bb";
      when "100111010" => romdata <= x"c9";
      when "100111011" => romdata <= x"58";
      when "100111100" => romdata <= x"2d";
      when "100111101" => romdata <= x"bc";
      when "100111110" => romdata <= x"ce";
      when "100111111" => romdata <= x"5f";
      when "101000000" => romdata <= x"70";
      when "101000001" => romdata <= x"e1";
      when "101000010" => romdata <= x"93";
      when "101000011" => romdata <= x"02";
      when "101000100" => romdata <= x"77";
      when "101000101" => romdata <= x"e6";
      when "101000110" => romdata <= x"94";
      when "101000111" => romdata <= x"05";
      when "101001000" => romdata <= x"7e";
      when "101001001" => romdata <= x"ef";
      when "101001010" => romdata <= x"9d";
      when "101001011" => romdata <= x"0c";
      when "101001100" => romdata <= x"79";
      when "101001101" => romdata <= x"e8";
      when "101001110" => romdata <= x"9a";
      when "101001111" => romdata <= x"0b";
      when "101010000" => romdata <= x"6c";
      when "101010001" => romdata <= x"fd";
      when "101010010" => romdata <= x"8f";
      when "101010011" => romdata <= x"1e";
      when "101010100" => romdata <= x"6b";
      when "101010101" => romdata <= x"fa";
      when "101010110" => romdata <= x"88";
      when "101010111" => romdata <= x"19";
      when "101011000" => romdata <= x"62";
      when "101011001" => romdata <= x"f3";
      when "101011010" => romdata <= x"81";
      when "101011011" => romdata <= x"10";
      when "101011100" => romdata <= x"65";
      when "101011101" => romdata <= x"f4";
      when "101011110" => romdata <= x"86";
      when "101011111" => romdata <= x"17";
      when "101100000" => romdata <= x"48";
      when "101100001" => romdata <= x"d9";
      when "101100010" => romdata <= x"ab";
      when "101100011" => romdata <= x"3a";
      when "101100100" => romdata <= x"4f";
      when "101100101" => romdata <= x"de";
      when "101100110" => romdata <= x"ac";
      when "101100111" => romdata <= x"3d";
      when "101101000" => romdata <= x"46";
      when "101101001" => romdata <= x"d7";
      when "101101010" => romdata <= x"a5";
      when "101101011" => romdata <= x"34";
      when "101101100" => romdata <= x"41";
      when "101101101" => romdata <= x"d0";
      when "101101110" => romdata <= x"a2";
      when "101101111" => romdata <= x"33";
      when "101110000" => romdata <= x"54";
      when "101110001" => romdata <= x"c5";
      when "101110010" => romdata <= x"b7";
      when "101110011" => romdata <= x"26";
      when "101110100" => romdata <= x"53";
      when "101110101" => romdata <= x"c2";
      when "101110110" => romdata <= x"b0";
      when "101110111" => romdata <= x"21";
      when "101111000" => romdata <= x"5a";
      when "101111001" => romdata <= x"cb";
      when "101111010" => romdata <= x"b9";
      when "101111011" => romdata <= x"28";
      when "101111100" => romdata <= x"5d";
      when "101111101" => romdata <= x"cc";
      when "101111110" => romdata <= x"be";
      when "101111111" => romdata <= x"2f";
      when "110000000" => romdata <= x"e0";
      when "110000001" => romdata <= x"71";
      when "110000010" => romdata <= x"03";
      when "110000011" => romdata <= x"92";
      when "110000100" => romdata <= x"e7";
      when "110000101" => romdata <= x"76";
      when "110000110" => romdata <= x"04";
      when "110000111" => romdata <= x"95";
      when "110001000" => romdata <= x"ee";
      when "110001001" => romdata <= x"7f";
      when "110001010" => romdata <= x"0d";
      when "110001011" => romdata <= x"9c";
      when "110001100" => romdata <= x"e9";
      when "110001101" => romdata <= x"78";
      when "110001110" => romdata <= x"0a";
      when "110001111" => romdata <= x"9b";
      when "110010000" => romdata <= x"fc";
      when "110010001" => romdata <= x"6d";
      when "110010010" => romdata <= x"1f";
      when "110010011" => romdata <= x"8e";
      when "110010100" => romdata <= x"fb";
      when "110010101" => romdata <= x"6a";
      when "110010110" => romdata <= x"18";
      when "110010111" => romdata <= x"89";
      when "110011000" => romdata <= x"f2";
      when "110011001" => romdata <= x"63";
      when "110011010" => romdata <= x"11";
      when "110011011" => romdata <= x"80";
      when "110011100" => romdata <= x"f5";
      when "110011101" => romdata <= x"64";
      when "110011110" => romdata <= x"16";
      when "110011111" => romdata <= x"87";
      when "110100000" => romdata <= x"d8";
      when "110100001" => romdata <= x"49";
      when "110100010" => romdata <= x"3b";
      when "110100011" => romdata <= x"aa";
      when "110100100" => romdata <= x"df";
      when "110100101" => romdata <= x"4e";
      when "110100110" => romdata <= x"3c";
      when "110100111" => romdata <= x"ad";
      when "110101000" => romdata <= x"d6";
      when "110101001" => romdata <= x"47";
      when "110101010" => romdata <= x"35";
      when "110101011" => romdata <= x"a4";
      when "110101100" => romdata <= x"d1";
      when "110101101" => romdata <= x"40";
      when "110101110" => romdata <= x"32";
      when "110101111" => romdata <= x"a3";
      when "110110000" => romdata <= x"c4";
      when "110110001" => romdata <= x"55";
      when "110110010" => romdata <= x"27";
      when "110110011" => romdata <= x"b6";
      when "110110100" => romdata <= x"c3";
      when "110110101" => romdata <= x"52";
      when "110110110" => romdata <= x"20";
      when "110110111" => romdata <= x"b1";
      when "110111000" => romdata <= x"ca";
      when "110111001" => romdata <= x"5b";
      when "110111010" => romdata <= x"29";
      when "110111011" => romdata <= x"b8";
      when "110111100" => romdata <= x"cd";
      when "110111101" => romdata <= x"5c";
      when "110111110" => romdata <= x"2e";
      when "110111111" => romdata <= x"bf";
      when "111000000" => romdata <= x"90";
      when "111000001" => romdata <= x"01";
      when "111000010" => romdata <= x"73";
      when "111000011" => romdata <= x"e2";
      when "111000100" => romdata <= x"97";
      when "111000101" => romdata <= x"06";
      when "111000110" => romdata <= x"74";
      when "111000111" => romdata <= x"e5";
      when "111001000" => romdata <= x"9e";
      when "111001001" => romdata <= x"0f";
      when "111001010" => romdata <= x"7d";
      when "111001011" => romdata <= x"ec";
      when "111001100" => romdata <= x"99";
      when "111001101" => romdata <= x"08";
      when "111001110" => romdata <= x"7a";
      when "111001111" => romdata <= x"eb";
      when "111010000" => romdata <= x"8c";
      when "111010001" => romdata <= x"1d";
      when "111010010" => romdata <= x"6f";
      when "111010011" => romdata <= x"fe";
      when "111010100" => romdata <= x"8b";
      when "111010101" => romdata <= x"1a";
      when "111010110" => romdata <= x"68";
      when "111010111" => romdata <= x"f9";
      when "111011000" => romdata <= x"82";
      when "111011001" => romdata <= x"13";
      when "111011010" => romdata <= x"61";
      when "111011011" => romdata <= x"f0";
      when "111011100" => romdata <= x"85";
      when "111011101" => romdata <= x"14";
      when "111011110" => romdata <= x"66";
      when "111011111" => romdata <= x"f7";
      when "111100000" => romdata <= x"a8";
      when "111100001" => romdata <= x"39";
      when "111100010" => romdata <= x"4b";
      when "111100011" => romdata <= x"da";
      when "111100100" => romdata <= x"af";
      when "111100101" => romdata <= x"3e";
      when "111100110" => romdata <= x"4c";
      when "111100111" => romdata <= x"dd";
      when "111101000" => romdata <= x"a6";
      when "111101001" => romdata <= x"37";
      when "111101010" => romdata <= x"45";
      when "111101011" => romdata <= x"d4";
      when "111101100" => romdata <= x"a1";
      when "111101101" => romdata <= x"30";
      when "111101110" => romdata <= x"42";
      when "111101111" => romdata <= x"d3";
      when "111110000" => romdata <= x"b4";
      when "111110001" => romdata <= x"25";
      when "111110010" => romdata <= x"57";
      when "111110011" => romdata <= x"c6";
      when "111110100" => romdata <= x"b3";
      when "111110101" => romdata <= x"22";
      when "111110110" => romdata <= x"50";
      when "111110111" => romdata <= x"c1";
      when "111111000" => romdata <= x"ba";
      when "111111001" => romdata <= x"2b";
      when "111111010" => romdata <= x"59";
      when "111111011" => romdata <= x"c8";
      when "111111100" => romdata <= x"bd";
      when "111111101" => romdata <= x"2c";
      when "111111110" => romdata <= x"5e";
      when "111111111" => romdata <= x"cf";
      when others      => romdata <= (others => '-');
    end case;
  end process comb;

  seq: process (clock) is
  begin  -- process seq
    if rising_edge(clock) then
      readData <= romdata;
    end if;
  end process seq;

end architecture rtl;

//--------------------------------------------------------------------
//
//  Description:  Cell Verilog models for mk180rtsc
//  Revision:     Rev: 1.02
//  Date:         Nov 30 2011
//
//--------------------------------------------------------------------

`timescale 1ns/10ps
`celldefine
module RT8_AA01D2 (Z, A1, A2, B, C);
input  A1 ;
input  A2 ;
input  B ;
input  C ;
output Z ;

   and (I0_out, A1, A2);
   or  (I1_out, I0_out, B);
   and (Z, I1_out, C);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$B$Z = 1.0,
       tphhl$B$Z = 1.0,
       tpllh$C$Z = 1.0,
       tphhl$C$Z = 1.0,
       tpllh$B$Z$A1_EQ_0_AN_A2_EQ_0_AN_C_EQ_1 = 1.0,
       tphhl$B$Z$A1_EQ_0_AN_A2_EQ_0_AN_C_EQ_1 = 1.0,
       tpllh$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_1 = 1.0,
       tphhl$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_1 = 1.0,
       tpllh$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_1 = 1.0,
       tphhl$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_1 = 1.0,
       tpllh$C$Z$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_1 = 1.0,
       tphhl$C$Z$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_1 = 1.0,
       tpllh$C$Z$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_1 = 1.0,
       tphhl$C$Z$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_1 = 1.0;

     // path delays


     if (A1 == 1'b1 && A2 == 1'b1 && B == 1'b1)
       (C *> Z) = (tpllh$C$Z$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_1, tphhl$C$Z$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b1)
       (C *> Z) = (tpllh$C$Z$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_1, tphhl$C$Z$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_1);
     ifnone
       (C *> Z) = (tpllh$C$Z,tphhl$C$Z);

     if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b1)
       (B *> Z) = (tpllh$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_1, tphhl$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b1)
       (B *> Z) = (tpllh$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_1, tphhl$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && C == 1'b1)
       (B *> Z) = (tpllh$B$Z$A1_EQ_0_AN_A2_EQ_0_AN_C_EQ_1, tphhl$B$Z$A1_EQ_0_AN_A2_EQ_0_AN_C_EQ_1);
     ifnone
       (B *> Z) = (tpllh$B$Z,tphhl$B$Z);

     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AA01D4 (Z, A1, A2, B, C);
input  A1 ;
input  A2 ;
input  B ;
input  C ;
output Z ;

   and (I0_out, A1, A2);
   or  (I1_out, I0_out, B);
   and (Z, I1_out, C);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$B$Z = 1.0,
       tphhl$B$Z = 1.0,
       tpllh$C$Z = 1.0,
       tphhl$C$Z = 1.0,
       tpllh$B$Z$A1_EQ_0_AN_A2_EQ_0_AN_C_EQ_1 = 1.0,
       tphhl$B$Z$A1_EQ_0_AN_A2_EQ_0_AN_C_EQ_1 = 1.0,
       tpllh$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_1 = 1.0,
       tphhl$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_1 = 1.0,
       tpllh$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_1 = 1.0,
       tphhl$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_1 = 1.0,
       tpllh$C$Z$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_1 = 1.0,
       tphhl$C$Z$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_1 = 1.0,
       tpllh$C$Z$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_1 = 1.0,
       tphhl$C$Z$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_1 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && B == 1'b1)
       (C *> Z) = (tpllh$C$Z$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_1, tphhl$C$Z$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b1)
       (C *> Z) = (tpllh$C$Z$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_1, tphhl$C$Z$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_1);
     ifnone
       (C *> Z) = (tpllh$C$Z,tphhl$C$Z);

     if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b1)
       (B *> Z) = (tpllh$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_1, tphhl$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b1)
       (B *> Z) = (tpllh$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_1, tphhl$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && C == 1'b1)
       (B *> Z) = (tpllh$B$Z$A1_EQ_0_AN_A2_EQ_0_AN_C_EQ_1, tphhl$B$Z$A1_EQ_0_AN_A2_EQ_0_AN_C_EQ_1);
     ifnone
       (B *> Z) = (tpllh$B$Z,tphhl$B$Z);

     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AAN1D1 (ZN, A1, A2, B, C);
input  A1 ;
input  A2 ;
input  B ;
input  C ;
output ZN ;

   and (I0_out, A1, A2);
   or  (I1_out, I0_out, B);
   and (I2_out, I1_out, C);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$B$ZN = 1.0,
       tphlh$B$ZN = 1.0,
       tplhl$C$ZN = 1.0,
       tphlh$C$ZN = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_C_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_C_EQ_1 = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_1 = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_1 = 1.0,
       tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_1 = 1.0,
       tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_1 = 1.0,
       tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_1 = 1.0,
       tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_1 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && B == 1'b1)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_1, tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b1)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_1, tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_1);
     ifnone
       (C *> ZN) = (tphlh$C$ZN,tplhl$C$ZN);

     if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_1, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_1, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && C == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_C_EQ_1, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_C_EQ_1);
     ifnone
       (B *> ZN) = (tphlh$B$ZN,tplhl$B$ZN);

     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AAN1D2 (ZN, A1, A2, B, C);
input  A1 ;
input  A2 ;
input  B ;
input  C ;
output ZN ;

   and (I0_out, A1, A2);
   or  (I1_out, I0_out, B);
   and (I2_out, I1_out, C);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$B$ZN = 1.0,
       tphlh$B$ZN = 1.0,
       tplhl$C$ZN = 1.0,
       tphlh$C$ZN = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_C_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_C_EQ_1 = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_1 = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_1 = 1.0,
       tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_1 = 1.0,
       tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_1 = 1.0,
       tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_1 = 1.0,
       tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_1 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && B == 1'b1)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_1, tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b1)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_1, tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_1);
     ifnone
       (C *> ZN) = (tphlh$C$ZN,tplhl$C$ZN);

     if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_1, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_1, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && C == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_C_EQ_1, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_C_EQ_1);
     ifnone
       (B *> ZN) = (tphlh$B$ZN,tplhl$B$ZN);

     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AAN1D4 (ZN, A1, A2, B, C);
input  A1 ;
input  A2 ;
input  B ;
input  C ;
output ZN ;

   and (I0_out, A1, A2);
   or  (I1_out, I0_out, B);
   and (I2_out, I1_out, C);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$B$ZN = 1.0,
       tphlh$B$ZN = 1.0,
       tplhl$C$ZN = 1.0,
       tphlh$C$ZN = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_C_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_C_EQ_1 = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_1 = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_1 = 1.0,
       tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_1 = 1.0,
       tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_1 = 1.0,
       tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_1 = 1.0,
       tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_1 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && B == 1'b1)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_1, tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b1)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_1, tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_1);
     ifnone
       (C *> ZN) = (tphlh$C$ZN,tplhl$C$ZN);

     if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_1, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_1, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && C == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_C_EQ_1, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_C_EQ_1);
     ifnone
       (B *> ZN) = (tphlh$B$ZN,tplhl$B$ZN);

     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AN02D1 (Z, A1, A2);
input  A1 ;
input  A2 ;
output Z ;

   and (Z, A1, A2);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0;

     // path delays
     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AN02D2 (Z, A1, A2);
input  A1 ;
input  A2 ;
output Z ;

   and (Z, A1, A2);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0;

     // path delays
     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AN02D4 (Z, A1, A2);
input  A1 ;
input  A2 ;
output Z ;

   and (Z, A1, A2);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0;

     // path delays
     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AN03D1 (Z, A1, A2, A3);
input  A1 ;
input  A2 ;
input  A3 ;
output Z ;

   and (Z, A1, A2, A3);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$A3$Z = 1.0,
       tphhl$A3$Z = 1.0;

     // path delays
     (A3 *> Z) = (tpllh$A3$Z, tphhl$A3$Z);
     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AN03D2 (Z, A1, A2, A3);
input  A1 ;
input  A2 ;
input  A3 ;
output Z ;

   and (Z, A1, A2, A3);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$A3$Z = 1.0,
       tphhl$A3$Z = 1.0;

     // path delays
     (A3 *> Z) = (tpllh$A3$Z, tphhl$A3$Z);
     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AN03D4 (Z, A1, A2, A3);
input  A1 ;
input  A2 ;
input  A3 ;
output Z ;

   and (Z, A1, A2, A3);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$A3$Z = 1.0,
       tphhl$A3$Z = 1.0;

     // path delays
     (A3 *> Z) = (tpllh$A3$Z, tphhl$A3$Z);
     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AN04D1 (Z, A1, A2, A3, A4);
input  A1 ;
input  A2 ;
input  A3 ;
input  A4 ;
output Z ;

   and (Z, A1, A2, A3, A4);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$A3$Z = 1.0,
       tphhl$A3$Z = 1.0,
       tpllh$A4$Z = 1.0,
       tphhl$A4$Z = 1.0;

     // path delays
     (A4 *> Z) = (tpllh$A4$Z, tphhl$A4$Z);
     (A3 *> Z) = (tpllh$A3$Z, tphhl$A3$Z);
     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AN04D2 (Z, A1, A2, A3, A4);
input  A1 ;
input  A2 ;
input  A3 ;
input  A4 ;
output Z ;

   and (Z, A1, A2, A3, A4);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$A3$Z = 1.0,
       tphhl$A3$Z = 1.0,
       tpllh$A4$Z = 1.0,
       tphhl$A4$Z = 1.0;

     // path delays
     (A4 *> Z) = (tpllh$A4$Z, tphhl$A4$Z);
     (A3 *> Z) = (tpllh$A3$Z, tphhl$A3$Z);
     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AN04D4 (Z, A1, A2, A3, A4);
input  A1 ;
input  A2 ;
input  A3 ;
input  A4 ;
output Z ;

   and (Z, A1, A2, A3, A4);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$A3$Z = 1.0,
       tphhl$A3$Z = 1.0,
       tpllh$A4$Z = 1.0,
       tphhl$A4$Z = 1.0;

     // path delays
     (A4 *> Z) = (tpllh$A4$Z, tphhl$A4$Z);
     (A3 *> Z) = (tpllh$A3$Z, tphhl$A3$Z);
     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AN06D2 (Z, A1, A2, A3, A4, A5, A6);
input  A1 ;
input  A2 ;
input  A3 ;
input  A4 ;
input  A5 ;
input  A6 ;
output Z ;

   and (Z, A1, A2, A3, A4, A5, A6);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$A3$Z = 1.0,
       tphhl$A3$Z = 1.0,
       tpllh$A4$Z = 1.0,
       tphhl$A4$Z = 1.0,
       tpllh$A5$Z = 1.0,
       tphhl$A5$Z = 1.0,
       tpllh$A6$Z = 1.0,
       tphhl$A6$Z = 1.0;

     // path delays
     (A6 *> Z) = (tpllh$A6$Z, tphhl$A6$Z);
     (A5 *> Z) = (tpllh$A5$Z, tphhl$A5$Z);
     (A4 *> Z) = (tpllh$A4$Z, tphhl$A4$Z);
     (A3 *> Z) = (tpllh$A3$Z, tphhl$A3$Z);
     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AN06D4 (Z, A1, A2, A3, A4, A5, A6);
input  A1 ;
input  A2 ;
input  A3 ;
input  A4 ;
input  A5 ;
input  A6 ;
output Z ;

   and (Z, A1, A2, A3, A4, A5, A6);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$A3$Z = 1.0,
       tphhl$A3$Z = 1.0,
       tpllh$A4$Z = 1.0,
       tphhl$A4$Z = 1.0,
       tpllh$A5$Z = 1.0,
       tphhl$A5$Z = 1.0,
       tpllh$A6$Z = 1.0,
       tphhl$A6$Z = 1.0;

     // path delays
     (A6 *> Z) = (tpllh$A6$Z, tphhl$A6$Z);
     (A5 *> Z) = (tpllh$A5$Z, tphhl$A5$Z);
     (A4 *> Z) = (tpllh$A4$Z, tphhl$A4$Z);
     (A3 *> Z) = (tpllh$A3$Z, tphhl$A3$Z);
     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AN08D2 (Z, A1, A2, A3, A4, A5, A6, A7, A8);
input  A1 ;
input  A2 ;
input  A3 ;
input  A4 ;
input  A5 ;
input  A6 ;
input  A7 ;
input  A8 ;
output Z ;

   and (Z, A1, A2, A3, A4, A5, A6, A7, A8);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$A3$Z = 1.0,
       tphhl$A3$Z = 1.0,
       tpllh$A4$Z = 1.0,
       tphhl$A4$Z = 1.0,
       tpllh$A5$Z = 1.0,
       tphhl$A5$Z = 1.0,
       tpllh$A6$Z = 1.0,
       tphhl$A6$Z = 1.0,
       tpllh$A7$Z = 1.0,
       tphhl$A7$Z = 1.0,
       tpllh$A8$Z = 1.0,
       tphhl$A8$Z = 1.0;

     // path delays
     (A8 *> Z) = (tpllh$A8$Z, tphhl$A8$Z);
     (A7 *> Z) = (tpllh$A7$Z, tphhl$A7$Z);
     (A6 *> Z) = (tpllh$A6$Z, tphhl$A6$Z);
     (A5 *> Z) = (tpllh$A5$Z, tphhl$A5$Z);
     (A4 *> Z) = (tpllh$A4$Z, tphhl$A4$Z);
     (A3 *> Z) = (tpllh$A3$Z, tphhl$A3$Z);
     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AN08D4 (Z, A1, A2, A3, A4, A5, A6, A7, A8);
input  A1 ;
input  A2 ;
input  A3 ;
input  A4 ;
input  A5 ;
input  A6 ;
input  A7 ;
input  A8 ;
output Z ;

   and (Z, A1, A2, A3, A4, A5, A6, A7, A8);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$A3$Z = 1.0,
       tphhl$A3$Z = 1.0,
       tpllh$A4$Z = 1.0,
       tphhl$A4$Z = 1.0,
       tpllh$A5$Z = 1.0,
       tphhl$A5$Z = 1.0,
       tpllh$A6$Z = 1.0,
       tphhl$A6$Z = 1.0,
       tpllh$A7$Z = 1.0,
       tphhl$A7$Z = 1.0,
       tpllh$A8$Z = 1.0,
       tphhl$A8$Z = 1.0;

     // path delays
     (A8 *> Z) = (tpllh$A8$Z, tphhl$A8$Z);
     (A7 *> Z) = (tpllh$A7$Z, tphhl$A7$Z);
     (A6 *> Z) = (tpllh$A6$Z, tphhl$A6$Z);
     (A5 *> Z) = (tpllh$A5$Z, tphhl$A5$Z);
     (A4 *> Z) = (tpllh$A4$Z, tphhl$A4$Z);
     (A3 *> Z) = (tpllh$A3$Z, tphhl$A3$Z);
     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AO01D2 (Z, A1, A2, B);
input  A1 ;
input  A2 ;
input  B ;
output Z ;

   and (I0_out, A1, A2);
   or  (Z, I0_out, B);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$B$Z = 1.0,
       tphhl$B$Z = 1.0,
       tpllh$B$Z$A1_EQ_0_AN_A2_EQ_0 = 1.0,
       tphhl$B$Z$A1_EQ_0_AN_A2_EQ_0 = 1.0,
       tpllh$B$Z$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tphhl$B$Z$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tpllh$B$Z$A1_EQ_1_AN_A2_EQ_0 = 1.0,
       tphhl$B$Z$A1_EQ_1_AN_A2_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b0)
       (B *> Z) = (tpllh$B$Z$A1_EQ_1_AN_A2_EQ_0, tphhl$B$Z$A1_EQ_1_AN_A2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1)
       (B *> Z) = (tpllh$B$Z$A1_EQ_0_AN_A2_EQ_1, tphhl$B$Z$A1_EQ_0_AN_A2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0)
       (B *> Z) = (tpllh$B$Z$A1_EQ_0_AN_A2_EQ_0, tphhl$B$Z$A1_EQ_0_AN_A2_EQ_0);
     ifnone
       (B *> Z) = (tpllh$B$Z,tphhl$B$Z);

     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AO01D4 (Z, A1, A2, B);
input  A1 ;
input  A2 ;
input  B ;
output Z ;

   and (I0_out, A1, A2);
   or  (Z, I0_out, B);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$B$Z = 1.0,
       tphhl$B$Z = 1.0,
       tpllh$B$Z$A1_EQ_0_AN_A2_EQ_0 = 1.0,
       tphhl$B$Z$A1_EQ_0_AN_A2_EQ_0 = 1.0,
       tpllh$B$Z$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tphhl$B$Z$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tpllh$B$Z$A1_EQ_1_AN_A2_EQ_0 = 1.0,
       tphhl$B$Z$A1_EQ_1_AN_A2_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b0)
       (B *> Z) = (tpllh$B$Z$A1_EQ_1_AN_A2_EQ_0, tphhl$B$Z$A1_EQ_1_AN_A2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1)
       (B *> Z) = (tpllh$B$Z$A1_EQ_0_AN_A2_EQ_1, tphhl$B$Z$A1_EQ_0_AN_A2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0)
       (B *> Z) = (tpllh$B$Z$A1_EQ_0_AN_A2_EQ_0, tphhl$B$Z$A1_EQ_0_AN_A2_EQ_0);
     ifnone
       (B *> Z) = (tpllh$B$Z,tphhl$B$Z);

     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AO02D2 (Z, A1, A2, B1, B2);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
output Z ;

   and (I0_out, A1, A2);
   and (I1_out, B1, B2);
   or  (Z, I0_out, I1_out);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$B1$Z = 1.0,
       tphhl$B1$Z = 1.0,
       tpllh$B2$Z = 1.0,
       tphhl$B2$Z = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1);
     ifnone
       (B2 *> Z) = (tpllh$B2$Z,tphhl$B2$Z);

     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1);
     ifnone
       (B1 *> Z) = (tpllh$B1$Z,tphhl$B1$Z);

     if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A2 *> Z) = (tpllh$A2$Z,tphhl$A2$Z);

     if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A1 *> Z) = (tpllh$A1$Z,tphhl$A1$Z);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AO02D4 (Z, A1, A2, B1, B2);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
output Z ;

   and (I0_out, A1, A2);
   and (I1_out, B1, B2);
   or  (Z, I0_out, I1_out);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$B1$Z = 1.0,
       tphhl$B1$Z = 1.0,
       tpllh$B2$Z = 1.0,
       tphhl$B2$Z = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1);
     ifnone
       (B2 *> Z) = (tpllh$B2$Z,tphhl$B2$Z);

     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1);
     ifnone
       (B1 *> Z) = (tpllh$B1$Z,tphhl$B1$Z);

     if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A2 *> Z) = (tpllh$A2$Z,tphhl$A2$Z);

     if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A1 *> Z) = (tpllh$A1$Z,tphhl$A1$Z);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AO03D2 (Z, A1, A2, A3, B);
input  A1 ;
input  A2 ;
input  A3 ;
input  B ;
output Z ;

   and (I1_out, A1, A2, A3);
   or  (Z, I1_out, B);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$A3$Z = 1.0,
       tphhl$A3$Z = 1.0,
       tpllh$B$Z = 1.0,
       tphhl$B$Z = 1.0,
       tpllh$B$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0 = 1.0,
       tphhl$B$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0 = 1.0,
       tpllh$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1 = 1.0,
       tphhl$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1 = 1.0,
       tpllh$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1 = 1.0,
       tphhl$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1 = 1.0,
       tpllh$B$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0 = 1.0,
       tphhl$B$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
       (B *> Z) = (tpllh$B$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0, tphhl$B$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
       (B *> Z) = (tpllh$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1, tphhl$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
       (B *> Z) = (tpllh$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1, tphhl$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
       (B *> Z) = (tpllh$B$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0, tphhl$B$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0);
     ifnone
       (B *> Z) = (tpllh$B$Z,tphhl$B$Z);

     (A3 *> Z) = (tpllh$A3$Z, tphhl$A3$Z);
     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AO03D4 (Z, A1, A2, A3, B);
input  A1 ;
input  A2 ;
input  A3 ;
input  B ;
output Z ;

   and (I1_out, A1, A2, A3);
   or  (Z, I1_out, B);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$A3$Z = 1.0,
       tphhl$A3$Z = 1.0,
       tpllh$B$Z = 1.0,
       tphhl$B$Z = 1.0,
       tpllh$B$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0 = 1.0,
       tphhl$B$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0 = 1.0,
       tpllh$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1 = 1.0,
       tphhl$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1 = 1.0,
       tpllh$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1 = 1.0,
       tphhl$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1 = 1.0,
       tpllh$B$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0 = 1.0,
       tphhl$B$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
       (B *> Z) = (tpllh$B$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0, tphhl$B$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
       (B *> Z) = (tpllh$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1, tphhl$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
       (B *> Z) = (tpllh$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1, tphhl$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
       (B *> Z) = (tpllh$B$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0, tphhl$B$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0);
     ifnone
       (B *> Z) = (tpllh$B$Z,tphhl$B$Z);

     (A3 *> Z) = (tpllh$A3$Z, tphhl$A3$Z);
     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AO04D2 (Z, A1, A2, A3, B1, B2);
input  A1 ;
input  A2 ;
input  A3 ;
input  B1 ;
input  B2 ;
output Z ;

   and (I1_out, A1, A2, A3);
   and (I2_out, B1, B2);
   or  (Z, I1_out, I2_out);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$A3$Z = 1.0,
       tphhl$A3$Z = 1.0,
       tpllh$B1$Z = 1.0,
       tphhl$B1$Z = 1.0,
       tpllh$B2$Z = 1.0,
       tphhl$B2$Z = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tpllh$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_1 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_1 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1);
     ifnone
       (B2 *> Z) = (tpllh$B2$Z,tphhl$B2$Z);

     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_1, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_1, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_1, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_1, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_1);
     ifnone
       (B1 *> Z) = (tpllh$B1$Z,tphhl$B1$Z);

     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A3 *> Z) = (tpllh$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A3 *> Z) = (tpllh$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (A3 *> Z) = (tpllh$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tphhl$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A3 *> Z) = (tpllh$A3$Z,tphhl$A3$Z);

     if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tphhl$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A2 *> Z) = (tpllh$A2$Z,tphhl$A2$Z);

     if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tphhl$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A1 *> Z) = (tpllh$A1$Z,tphhl$A1$Z);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AO04D4 (Z, A1, A2, A3, B1, B2);
input  A1 ;
input  A2 ;
input  A3 ;
input  B1 ;
input  B2 ;
output Z ;

   and (I1_out, A1, A2, A3);
   and (I2_out, B1, B2);
   or  (Z, I1_out, I2_out);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$A3$Z = 1.0,
       tphhl$A3$Z = 1.0,
       tpllh$B1$Z = 1.0,
       tphhl$B1$Z = 1.0,
       tpllh$B2$Z = 1.0,
       tphhl$B2$Z = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tpllh$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_1 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_1 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1);
     ifnone
       (B2 *> Z) = (tpllh$B2$Z,tphhl$B2$Z);

     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_1, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_1, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_1, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_1, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_1);
     ifnone
       (B1 *> Z) = (tpllh$B1$Z,tphhl$B1$Z);

     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A3 *> Z) = (tpllh$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A3 *> Z) = (tpllh$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (A3 *> Z) = (tpllh$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tphhl$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A3 *> Z) = (tpllh$A3$Z,tphhl$A3$Z);

     if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tphhl$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A2 *> Z) = (tpllh$A2$Z,tphhl$A2$Z);

     if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tphhl$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A1 *> Z) = (tpllh$A1$Z,tphhl$A1$Z);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AO05D2 (Z, A1, A2, A3, B1, B2, B3);
input  A1 ;
input  A2 ;
input  A3 ;
input  B1 ;
input  B2 ;
input  B3 ;
output Z ;

   and (I1_out, A1, A2, A3);
   and (I3_out, B1, B2, B3);
   or  (Z, I1_out, I3_out);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$A3$Z = 1.0,
       tphhl$A3$Z = 1.0,
       tpllh$B1$Z = 1.0,
       tphhl$B1$Z = 1.0,
       tpllh$B2$Z = 1.0,
       tphhl$B2$Z = 1.0,
       tpllh$B3$Z = 1.0,
       tphhl$B3$Z = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tpllh$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphhl$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tpllh$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphhl$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tpllh$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tphhl$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tpllh$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tphhl$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B3_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B3_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B3_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B3_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1_AN_B3_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1_AN_B3_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1_AN_B3_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1_AN_B3_EQ_1 = 1.0,
       tpllh$B3$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$B3$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tpllh$B3$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$B3$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tpllh$B3$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$B3$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tpllh$B3$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$B3$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (B3 *> Z) = (tpllh$B3$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tphhl$B3$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
       (B3 *> Z) = (tpllh$B3$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1, tphhl$B3$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
       (B3 *> Z) = (tpllh$B3$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1, tphhl$B3$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (B3 *> Z) = (tpllh$B3$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tphhl$B3$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     ifnone
       (B3 *> Z) = (tpllh$B3$Z,tphhl$B3$Z);

     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1_AN_B3_EQ_1, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1_AN_B3_EQ_1, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B3_EQ_1, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B3_EQ_1, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B3_EQ_1);
     ifnone
       (B2 *> Z) = (tpllh$B2$Z,tphhl$B2$Z);

     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1);
     ifnone
       (B1 *> Z) = (tpllh$B1$Z,tphhl$B1$Z);

     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
       (A3 *> Z) = (tpllh$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0, tphhl$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
       (A3 *> Z) = (tpllh$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1, tphhl$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
       (A3 *> Z) = (tpllh$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1, tphhl$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
       (A3 *> Z) = (tpllh$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0, tphhl$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0);
     ifnone
       (A3 *> Z) = (tpllh$A3$Z,tphhl$A3$Z);

     if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0, tphhl$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0);
     if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1, tphhl$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1);
     if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1, tphhl$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0, tphhl$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0);
     ifnone
       (A2 *> Z) = (tpllh$A2$Z,tphhl$A2$Z);

     if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0, tphhl$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0);
     if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1, tphhl$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1);
     if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1, tphhl$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0, tphhl$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0);
     ifnone
       (A1 *> Z) = (tpllh$A1$Z,tphhl$A1$Z);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AO05D4 (Z, A1, A2, A3, B1, B2, B3);
input  A1 ;
input  A2 ;
input  A3 ;
input  B1 ;
input  B2 ;
input  B3 ;
output Z ;

   and (I1_out, A1, A2, A3);
   and (I3_out, B1, B2, B3);
   or  (Z, I1_out, I3_out);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$A3$Z = 1.0,
       tphhl$A3$Z = 1.0,
       tpllh$B1$Z = 1.0,
       tphhl$B1$Z = 1.0,
       tpllh$B2$Z = 1.0,
       tphhl$B2$Z = 1.0,
       tpllh$B3$Z = 1.0,
       tphhl$B3$Z = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tpllh$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphhl$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tpllh$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphhl$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tpllh$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tphhl$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tpllh$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tphhl$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B3_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B3_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B3_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B3_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1_AN_B3_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1_AN_B3_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1_AN_B3_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1_AN_B3_EQ_1 = 1.0,
       tpllh$B3$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$B3$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tpllh$B3$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$B3$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tpllh$B3$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$B3$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tpllh$B3$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$B3$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (B3 *> Z) = (tpllh$B3$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tphhl$B3$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
       (B3 *> Z) = (tpllh$B3$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1, tphhl$B3$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
       (B3 *> Z) = (tpllh$B3$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1, tphhl$B3$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (B3 *> Z) = (tpllh$B3$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tphhl$B3$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     ifnone
       (B3 *> Z) = (tpllh$B3$Z,tphhl$B3$Z);

     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1_AN_B3_EQ_1, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1_AN_B3_EQ_1, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B3_EQ_1, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B3_EQ_1, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B3_EQ_1);
     ifnone
       (B2 *> Z) = (tpllh$B2$Z,tphhl$B2$Z);

     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1);
     ifnone
       (B1 *> Z) = (tpllh$B1$Z,tphhl$B1$Z);

     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
       (A3 *> Z) = (tpllh$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0, tphhl$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
       (A3 *> Z) = (tpllh$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1, tphhl$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
       (A3 *> Z) = (tpllh$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1, tphhl$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
       (A3 *> Z) = (tpllh$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0, tphhl$A3$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0);
     ifnone
       (A3 *> Z) = (tpllh$A3$Z,tphhl$A3$Z);

     if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0, tphhl$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0);
     if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1, tphhl$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1);
     if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1, tphhl$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0, tphhl$A2$Z$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0);
     ifnone
       (A2 *> Z) = (tpllh$A2$Z,tphhl$A2$Z);

     if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0, tphhl$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0);
     if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1, tphhl$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1);
     if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1, tphhl$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0, tphhl$A1$Z$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0);
     ifnone
       (A1 *> Z) = (tpllh$A1$Z,tphhl$A1$Z);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AO06D2 (Z, A1, A2, B, C);
input  A1 ;
input  A2 ;
input  B ;
input  C ;
output Z ;

   and (I0_out, A1, A2);
   or  (Z, I0_out, B, C);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$B$Z = 1.0,
       tphhl$B$Z = 1.0,
       tpllh$C$Z = 1.0,
       tphhl$C$Z = 1.0,
       tpllh$B$Z$A1_EQ_0_AN_A2_EQ_0_AN_C_EQ_0 = 1.0,
       tphhl$B$Z$A1_EQ_0_AN_A2_EQ_0_AN_C_EQ_0 = 1.0,
       tpllh$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_0 = 1.0,
       tphhl$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_0 = 1.0,
       tpllh$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_0 = 1.0,
       tphhl$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_0 = 1.0,
       tpllh$C$Z$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_0 = 1.0,
       tphhl$C$Z$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_0 = 1.0,
       tpllh$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B_EQ_0 = 1.0,
       tphhl$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B_EQ_0 = 1.0,
       tpllh$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B_EQ_0 = 1.0,
       tphhl$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b0)
       (C *> Z) = (tpllh$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B_EQ_0, tphhl$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b0)
       (C *> Z) = (tpllh$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B_EQ_0, tphhl$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b0)
       (C *> Z) = (tpllh$C$Z$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_0, tphhl$C$Z$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_0);
     ifnone
       (C *> Z) = (tpllh$C$Z,tphhl$C$Z);

     if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b0)
       (B *> Z) = (tpllh$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_0, tphhl$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b0)
       (B *> Z) = (tpllh$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_0, tphhl$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && C == 1'b0)
       (B *> Z) = (tpllh$B$Z$A1_EQ_0_AN_A2_EQ_0_AN_C_EQ_0, tphhl$B$Z$A1_EQ_0_AN_A2_EQ_0_AN_C_EQ_0);
     ifnone
       (B *> Z) = (tpllh$B$Z,tphhl$B$Z);

     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AO06D4 (Z, A1, A2, B, C);
input  A1 ;
input  A2 ;
input  B ;
input  C ;
output Z ;

   and (I0_out, A1, A2);
   or  (Z, I0_out, B, C);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$B$Z = 1.0,
       tphhl$B$Z = 1.0,
       tpllh$C$Z = 1.0,
       tphhl$C$Z = 1.0,
       tpllh$B$Z$A1_EQ_0_AN_A2_EQ_0_AN_C_EQ_0 = 1.0,
       tphhl$B$Z$A1_EQ_0_AN_A2_EQ_0_AN_C_EQ_0 = 1.0,
       tpllh$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_0 = 1.0,
       tphhl$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_0 = 1.0,
       tpllh$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_0 = 1.0,
       tphhl$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_0 = 1.0,
       tpllh$C$Z$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_0 = 1.0,
       tphhl$C$Z$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_0 = 1.0,
       tpllh$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B_EQ_0 = 1.0,
       tphhl$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B_EQ_0 = 1.0,
       tpllh$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B_EQ_0 = 1.0,
       tphhl$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b0)
       (C *> Z) = (tpllh$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B_EQ_0, tphhl$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b0)
       (C *> Z) = (tpllh$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B_EQ_0, tphhl$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b0)
       (C *> Z) = (tpllh$C$Z$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_0, tphhl$C$Z$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_0);
     ifnone
       (C *> Z) = (tpllh$C$Z,tphhl$C$Z);

     if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b0)
       (B *> Z) = (tpllh$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_0, tphhl$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b0)
       (B *> Z) = (tpllh$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_0, tphhl$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && C == 1'b0)
       (B *> Z) = (tpllh$B$Z$A1_EQ_0_AN_A2_EQ_0_AN_C_EQ_0, tphhl$B$Z$A1_EQ_0_AN_A2_EQ_0_AN_C_EQ_0);
     ifnone
       (B *> Z) = (tpllh$B$Z,tphhl$B$Z);

     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AO07D2 (Z, A1, A2, B1, B2, C);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
input  C ;
output Z ;

   and (I0_out, A1, A2);
   and (I1_out, B1, B2);
   or  (Z, I0_out, I1_out, C);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$B1$Z = 1.0,
       tphhl$B1$Z = 1.0,
       tpllh$B2$Z = 1.0,
       tphhl$B2$Z = 1.0,
       tpllh$C$Z = 1.0,
       tphhl$C$Z = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C_EQ_0 = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_C_EQ_0 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_C_EQ_0 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C_EQ_0 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C_EQ_0 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C_EQ_0 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C_EQ_0 = 1.0,
       tpllh$C$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$C$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tpllh$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (C *> Z) = (tpllh$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (C *> Z) = (tpllh$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (C *> Z) = (tpllh$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (C *> Z) = (tpllh$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
       (C *> Z) = (tpllh$C$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0, tphhl$C$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (C *> Z) = (tpllh$C$Z,tphhl$C$Z);

     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C_EQ_0, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C == 1'b0)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C_EQ_0, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_C_EQ_0, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_C_EQ_0);
     ifnone
       (B2 *> Z) = (tpllh$B2$Z,tphhl$B2$Z);

     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C_EQ_0, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C == 1'b0)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C_EQ_0, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1_AN_C_EQ_0, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1_AN_C_EQ_0);
     ifnone
       (B1 *> Z) = (tpllh$B1$Z,tphhl$B1$Z);

     if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_0, tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_0);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_0, tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_0);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C_EQ_0, tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C_EQ_0);
     ifnone
       (A2 *> Z) = (tpllh$A2$Z,tphhl$A2$Z);

     if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_0, tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_0);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_0, tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_0);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C_EQ_0, tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C_EQ_0);
     ifnone
       (A1 *> Z) = (tpllh$A1$Z,tphhl$A1$Z);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AO07D4 (Z, A1, A2, B1, B2, C);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
input  C ;
output Z ;

   and (I0_out, A1, A2);
   and (I1_out, B1, B2);
   or  (Z, I0_out, I1_out, C);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$B1$Z = 1.0,
       tphhl$B1$Z = 1.0,
       tpllh$B2$Z = 1.0,
       tphhl$B2$Z = 1.0,
       tpllh$C$Z = 1.0,
       tphhl$C$Z = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C_EQ_0 = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_C_EQ_0 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_C_EQ_0 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C_EQ_0 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C_EQ_0 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C_EQ_0 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C_EQ_0 = 1.0,
       tpllh$C$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$C$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tpllh$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (C *> Z) = (tpllh$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (C *> Z) = (tpllh$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (C *> Z) = (tpllh$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (C *> Z) = (tpllh$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
       (C *> Z) = (tpllh$C$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0, tphhl$C$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (C *> Z) = (tpllh$C$Z,tphhl$C$Z);

     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C_EQ_0, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C == 1'b0)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C_EQ_0, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_C_EQ_0, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_C_EQ_0);
     ifnone
       (B2 *> Z) = (tpllh$B2$Z,tphhl$B2$Z);

     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C_EQ_0, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C == 1'b0)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C_EQ_0, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1_AN_C_EQ_0, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1_AN_C_EQ_0);
     ifnone
       (B1 *> Z) = (tpllh$B1$Z,tphhl$B1$Z);

     if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_0, tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_0);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_0, tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_0);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C_EQ_0, tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C_EQ_0);
     ifnone
       (A2 *> Z) = (tpllh$A2$Z,tphhl$A2$Z);

     if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_0, tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_0);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_0, tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_0);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C_EQ_0, tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C_EQ_0);
     ifnone
       (A1 *> Z) = (tpllh$A1$Z,tphhl$A1$Z);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AO08D2 (Z, A1, A2, B1, B2, C1, C2);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
input  C1 ;
input  C2 ;
output Z ;

   and (I0_out, C1, C2);
   and (I1_out, A1, A2);
   and (I3_out, B1, B2);
   or  (Z, I0_out, I1_out, I3_out);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$B1$Z = 1.0,
       tphhl$B1$Z = 1.0,
       tpllh$B2$Z = 1.0,
       tphhl$B2$Z = 1.0,
       tpllh$C1$Z = 1.0,
       tphhl$C1$Z = 1.0,
       tpllh$C2$Z = 1.0,
       tphhl$C2$Z = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_0 = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_0 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_0 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_0 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tpllh$C1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_C2_EQ_1 = 1.0,
       tphhl$C1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_C2_EQ_1 = 1.0,
       tpllh$C1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_1 = 1.0,
       tphhl$C1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_1 = 1.0,
       tpllh$C1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_1 = 1.0,
       tphhl$C1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_1 = 1.0,
       tpllh$C1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_1 = 1.0,
       tphhl$C1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_1 = 1.0,
       tpllh$C1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_1 = 1.0,
       tphhl$C1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_1 = 1.0,
       tpllh$C2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_1 = 1.0,
       tphhl$C2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_1 = 1.0,
       tpllh$C2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1 = 1.0,
       tphhl$C2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1 = 1.0,
       tpllh$C2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1 = 1.0,
       tphhl$C2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1 = 1.0,
       tpllh$C2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1 = 1.0,
       tphhl$C2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1 = 1.0,
       tpllh$C2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1 = 1.0,
       tphhl$C2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
       (C2 *> Z) = (tpllh$C2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1, tphhl$C2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
       (C2 *> Z) = (tpllh$C2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1, tphhl$C2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
       (C2 *> Z) = (tpllh$C2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1, tphhl$C2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
       (C2 *> Z) = (tpllh$C2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1, tphhl$C2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
       (C2 *> Z) = (tpllh$C2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_1, tphhl$C2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_1);
     ifnone
       (C2 *> Z) = (tpllh$C2$Z,tphhl$C2$Z);

     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
       (C1 *> Z) = (tpllh$C1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_1, tphhl$C1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
       (C1 *> Z) = (tpllh$C1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_1, tphhl$C1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
       (C1 *> Z) = (tpllh$C1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_1, tphhl$C1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
       (C1 *> Z) = (tpllh$C1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_1, tphhl$C1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
       (C1 *> Z) = (tpllh$C1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_C2_EQ_1, tphhl$C1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_C2_EQ_1);
     ifnone
       (C1 *> Z) = (tpllh$C1$Z,tphhl$C1$Z);

     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_0, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_0);
     ifnone
       (B2 *> Z) = (tpllh$B2$Z,tphhl$B2$Z);

     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_0, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_0);
     ifnone
       (B1 *> Z) = (tpllh$B1$Z,tphhl$B1$Z);

     if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0, tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1, tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0, tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1, tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_0, tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_0);
     ifnone
       (A2 *> Z) = (tpllh$A2$Z,tphhl$A2$Z);

     if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0, tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1, tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0, tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1, tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_0, tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_0);
     ifnone
       (A1 *> Z) = (tpllh$A1$Z,tphhl$A1$Z);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AO08D4 (Z, A1, A2, B1, B2, C1, C2);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
input  C1 ;
input  C2 ;
output Z ;

   and (I0_out, C1, C2);
   and (I1_out, A1, A2);
   and (I3_out, B1, B2);
   or  (Z, I0_out, I1_out, I3_out);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$B1$Z = 1.0,
       tphhl$B1$Z = 1.0,
       tpllh$B2$Z = 1.0,
       tphhl$B2$Z = 1.0,
       tpllh$C1$Z = 1.0,
       tphhl$C1$Z = 1.0,
       tpllh$C2$Z = 1.0,
       tphhl$C2$Z = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_0 = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_0 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_0 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_0 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tpllh$C1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_C2_EQ_1 = 1.0,
       tphhl$C1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_C2_EQ_1 = 1.0,
       tpllh$C1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_1 = 1.0,
       tphhl$C1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_1 = 1.0,
       tpllh$C1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_1 = 1.0,
       tphhl$C1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_1 = 1.0,
       tpllh$C1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_1 = 1.0,
       tphhl$C1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_1 = 1.0,
       tpllh$C1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_1 = 1.0,
       tphhl$C1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_1 = 1.0,
       tpllh$C2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_1 = 1.0,
       tphhl$C2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_1 = 1.0,
       tpllh$C2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1 = 1.0,
       tphhl$C2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1 = 1.0,
       tpllh$C2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1 = 1.0,
       tphhl$C2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1 = 1.0,
       tpllh$C2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1 = 1.0,
       tphhl$C2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1 = 1.0,
       tpllh$C2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1 = 1.0,
       tphhl$C2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
       (C2 *> Z) = (tpllh$C2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1, tphhl$C2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
       (C2 *> Z) = (tpllh$C2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1, tphhl$C2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
       (C2 *> Z) = (tpllh$C2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1, tphhl$C2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
       (C2 *> Z) = (tpllh$C2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1, tphhl$C2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
       (C2 *> Z) = (tpllh$C2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_1, tphhl$C2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_1);
     ifnone
       (C2 *> Z) = (tpllh$C2$Z,tphhl$C2$Z);

     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
       (C1 *> Z) = (tpllh$C1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_1, tphhl$C1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
       (C1 *> Z) = (tpllh$C1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_1, tphhl$C1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
       (C1 *> Z) = (tpllh$C1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_1, tphhl$C1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
       (C1 *> Z) = (tpllh$C1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_1, tphhl$C1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
       (C1 *> Z) = (tpllh$C1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_C2_EQ_1, tphhl$C1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_C2_EQ_1);
     ifnone
       (C1 *> Z) = (tpllh$C1$Z,tphhl$C1$Z);

     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_0, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_0);
     ifnone
       (B2 *> Z) = (tpllh$B2$Z,tphhl$B2$Z);

     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_0, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_0);
     ifnone
       (B1 *> Z) = (tpllh$B1$Z,tphhl$B1$Z);

     if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0, tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1, tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0, tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1, tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_0, tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_0);
     ifnone
       (A2 *> Z) = (tpllh$A2$Z,tphhl$A2$Z);

     if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0, tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1, tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0, tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1, tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_0, tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_0);
     ifnone
       (A1 *> Z) = (tpllh$A1$Z,tphhl$A1$Z);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AON1BBD1 (ZN, A1N, A2N, B);
input  A1N ;
input  A2N ;
input  B ;
output ZN ;

   or  (I0_out, A1N, A2N);
   not (I1_out, I0_out);
   or  (I2_out, I1_out, B);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tpllh$A1N$ZN = 1.0,
       tphhl$A1N$ZN = 1.0,
       tpllh$A2N$ZN = 1.0,
       tphhl$A2N$ZN = 1.0,
       tplhl$B$ZN = 1.0,
       tphlh$B$ZN = 1.0,
       tplhl$B$ZN$A1N_EQ_1_AN_A2N_EQ_1 = 1.0,
       tphlh$B$ZN$A1N_EQ_1_AN_A2N_EQ_1 = 1.0,
       tplhl$B$ZN$A1N_EQ_1_AN_A2N_EQ_0 = 1.0,
       tphlh$B$ZN$A1N_EQ_1_AN_A2N_EQ_0 = 1.0,
       tplhl$B$ZN$A1N_EQ_0_AN_A2N_EQ_1 = 1.0,
       tphlh$B$ZN$A1N_EQ_0_AN_A2N_EQ_1 = 1.0;

     // path delays
     if (A1N == 1'b1 && A2N == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1N_EQ_1_AN_A2N_EQ_1, tplhl$B$ZN$A1N_EQ_1_AN_A2N_EQ_1);
     if (A1N == 1'b1 && A2N == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1N_EQ_1_AN_A2N_EQ_0, tplhl$B$ZN$A1N_EQ_1_AN_A2N_EQ_0);
     if (A1N == 1'b0 && A2N == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1N_EQ_0_AN_A2N_EQ_1, tplhl$B$ZN$A1N_EQ_0_AN_A2N_EQ_1);
     ifnone
       (B *> ZN) = (tphlh$B$ZN,tplhl$B$ZN);

     (A2N *> ZN) = (tpllh$A2N$ZN, tphhl$A2N$ZN);
     (A1N *> ZN) = (tpllh$A1N$ZN, tphhl$A1N$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AON1BBD2 (ZN, A1N, A2N, B);
input  A1N ;
input  A2N ;
input  B ;
output ZN ;

   or  (I0_out, A1N, A2N);
   not (I1_out, I0_out);
   or  (I2_out, I1_out, B);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tpllh$A1N$ZN = 1.0,
       tphhl$A1N$ZN = 1.0,
       tpllh$A2N$ZN = 1.0,
       tphhl$A2N$ZN = 1.0,
       tplhl$B$ZN = 1.0,
       tphlh$B$ZN = 1.0,
       tplhl$B$ZN$A1N_EQ_1_AN_A2N_EQ_1 = 1.0,
       tphlh$B$ZN$A1N_EQ_1_AN_A2N_EQ_1 = 1.0,
       tplhl$B$ZN$A1N_EQ_1_AN_A2N_EQ_0 = 1.0,
       tphlh$B$ZN$A1N_EQ_1_AN_A2N_EQ_0 = 1.0,
       tplhl$B$ZN$A1N_EQ_0_AN_A2N_EQ_1 = 1.0,
       tphlh$B$ZN$A1N_EQ_0_AN_A2N_EQ_1 = 1.0;

     // path delays
     if (A1N == 1'b1 && A2N == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1N_EQ_1_AN_A2N_EQ_1, tplhl$B$ZN$A1N_EQ_1_AN_A2N_EQ_1);
     if (A1N == 1'b1 && A2N == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1N_EQ_1_AN_A2N_EQ_0, tplhl$B$ZN$A1N_EQ_1_AN_A2N_EQ_0);
     if (A1N == 1'b0 && A2N == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1N_EQ_0_AN_A2N_EQ_1, tplhl$B$ZN$A1N_EQ_0_AN_A2N_EQ_1);
     ifnone
       (B *> ZN) = (tphlh$B$ZN,tplhl$B$ZN);

     (A2N *> ZN) = (tpllh$A2N$ZN, tphhl$A2N$ZN);
     (A1N *> ZN) = (tpllh$A1N$ZN, tphhl$A1N$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AON1BBD4 (ZN, A1N, A2N, B);
input  A1N ;
input  A2N ;
input  B ;
output ZN ;

   or  (I0_out, A1N, A2N);
   not (I1_out, I0_out);
   or  (I2_out, I1_out, B);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tpllh$A1N$ZN = 1.0,
       tphhl$A1N$ZN = 1.0,
       tpllh$A2N$ZN = 1.0,
       tphhl$A2N$ZN = 1.0,
       tplhl$B$ZN = 1.0,
       tphlh$B$ZN = 1.0,
       tplhl$B$ZN$A1N_EQ_1_AN_A2N_EQ_1 = 1.0,
       tphlh$B$ZN$A1N_EQ_1_AN_A2N_EQ_1 = 1.0,
       tplhl$B$ZN$A1N_EQ_1_AN_A2N_EQ_0 = 1.0,
       tphlh$B$ZN$A1N_EQ_1_AN_A2N_EQ_0 = 1.0,
       tplhl$B$ZN$A1N_EQ_0_AN_A2N_EQ_1 = 1.0,
       tphlh$B$ZN$A1N_EQ_0_AN_A2N_EQ_1 = 1.0;

     // path delays
     if (A1N == 1'b1 && A2N == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1N_EQ_1_AN_A2N_EQ_1, tplhl$B$ZN$A1N_EQ_1_AN_A2N_EQ_1);
     if (A1N == 1'b1 && A2N == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1N_EQ_1_AN_A2N_EQ_0, tplhl$B$ZN$A1N_EQ_1_AN_A2N_EQ_0);
     if (A1N == 1'b0 && A2N == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1N_EQ_0_AN_A2N_EQ_1, tplhl$B$ZN$A1N_EQ_0_AN_A2N_EQ_1);
     ifnone
       (B *> ZN) = (tphlh$B$ZN,tplhl$B$ZN);

     (A2N *> ZN) = (tpllh$A2N$ZN, tphhl$A2N$ZN);
     (A1N *> ZN) = (tpllh$A1N$ZN, tphhl$A1N$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AON1BD1 (ZN, A1, A2, BN);
input  A1 ;
input  A2 ;
input  BN ;
output ZN ;

   and (I0_out, A1, A2);
   not (I1_out, I0_out);
   and (ZN, I1_out, BN);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tpllh$BN$ZN = 1.0,
       tphhl$BN$ZN = 1.0,
       tpllh$BN$ZN$A1_EQ_0_AN_A2_EQ_0 = 1.0,
       tphhl$BN$ZN$A1_EQ_0_AN_A2_EQ_0 = 1.0,
       tpllh$BN$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tphhl$BN$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tpllh$BN$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0,
       tphhl$BN$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b0)
       (BN *> ZN) = (tpllh$BN$ZN$A1_EQ_1_AN_A2_EQ_0, tphhl$BN$ZN$A1_EQ_1_AN_A2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1)
       (BN *> ZN) = (tpllh$BN$ZN$A1_EQ_0_AN_A2_EQ_1, tphhl$BN$ZN$A1_EQ_0_AN_A2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0)
       (BN *> ZN) = (tpllh$BN$ZN$A1_EQ_0_AN_A2_EQ_0, tphhl$BN$ZN$A1_EQ_0_AN_A2_EQ_0);
     ifnone
       (BN *> ZN) = (tpllh$BN$ZN,tphhl$BN$ZN);

     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AON1BD2 (ZN, A1, A2, BN);
input  A1 ;
input  A2 ;
input  BN ;
output ZN ;

   and (I0_out, A1, A2);
   not (I1_out, I0_out);
   and (ZN, I1_out, BN);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tpllh$BN$ZN = 1.0,
       tphhl$BN$ZN = 1.0,
       tpllh$BN$ZN$A1_EQ_0_AN_A2_EQ_0 = 1.0,
       tphhl$BN$ZN$A1_EQ_0_AN_A2_EQ_0 = 1.0,
       tpllh$BN$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tphhl$BN$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tpllh$BN$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0,
       tphhl$BN$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b0)
       (BN *> ZN) = (tpllh$BN$ZN$A1_EQ_1_AN_A2_EQ_0, tphhl$BN$ZN$A1_EQ_1_AN_A2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1)
       (BN *> ZN) = (tpllh$BN$ZN$A1_EQ_0_AN_A2_EQ_1, tphhl$BN$ZN$A1_EQ_0_AN_A2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0)
       (BN *> ZN) = (tpllh$BN$ZN$A1_EQ_0_AN_A2_EQ_0, tphhl$BN$ZN$A1_EQ_0_AN_A2_EQ_0);
     ifnone
       (BN *> ZN) = (tpllh$BN$ZN,tphhl$BN$ZN);

     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AON1BD4 (ZN, A1, A2, BN);
input  A1 ;
input  A2 ;
input  BN ;
output ZN ;

   and (I0_out, A1, A2);
   not (I1_out, I0_out);
   and (ZN, I1_out, BN);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tpllh$BN$ZN = 1.0,
       tphhl$BN$ZN = 1.0,
       tpllh$BN$ZN$A1_EQ_0_AN_A2_EQ_0 = 1.0,
       tphhl$BN$ZN$A1_EQ_0_AN_A2_EQ_0 = 1.0,
       tpllh$BN$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tphhl$BN$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tpllh$BN$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0,
       tphhl$BN$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b0)
       (BN *> ZN) = (tpllh$BN$ZN$A1_EQ_1_AN_A2_EQ_0, tphhl$BN$ZN$A1_EQ_1_AN_A2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1)
       (BN *> ZN) = (tpllh$BN$ZN$A1_EQ_0_AN_A2_EQ_1, tphhl$BN$ZN$A1_EQ_0_AN_A2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0)
       (BN *> ZN) = (tpllh$BN$ZN$A1_EQ_0_AN_A2_EQ_0, tphhl$BN$ZN$A1_EQ_0_AN_A2_EQ_0);
     ifnone
       (BN *> ZN) = (tpllh$BN$ZN,tphhl$BN$ZN);

     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AON1D1 (ZN, A1, A2, B);
input  A1 ;
input  A2 ;
input  B ;
output ZN ;

   and (I0_out, A1, A2);
   or  (I1_out, I0_out, B);
   not (ZN, I1_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$B$ZN = 1.0,
       tphlh$B$ZN = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_0 = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_0, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_0);
     ifnone
       (B *> ZN) = (tphlh$B$ZN,tplhl$B$ZN);

     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AON1D2 (ZN, A1, A2, B);
input  A1 ;
input  A2 ;
input  B ;
output ZN ;

   and (I0_out, A1, A2);
   or  (I1_out, I0_out, B);
   not (ZN, I1_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$B$ZN = 1.0,
       tphlh$B$ZN = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_0 = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_0, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_0);
     ifnone
       (B *> ZN) = (tphlh$B$ZN,tplhl$B$ZN);

     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AON1D4 (ZN, A1, A2, B);
input  A1 ;
input  A2 ;
input  B ;
output ZN ;

   and (I0_out, A1, A2);
   or  (I1_out, I0_out, B);
   not (ZN, I1_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$B$ZN = 1.0,
       tphlh$B$ZN = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_0 = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_0, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_0);
     ifnone
       (B *> ZN) = (tphlh$B$ZN,tplhl$B$ZN);

     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AON2BBD1 (ZN, A1N, A2N, B1, B2);
input  A1N ;
input  A2N ;
input  B1 ;
input  B2 ;
output ZN ;

   or  (I0_out, A1N, A2N);
   not (I1_out, I0_out);
   and (I2_out, B1, B2);
   or  (I3_out, I1_out, I2_out);
   not (ZN, I3_out);

   specify
     // delay parameters
     specparam
       tpllh$A1N$ZN = 1.0,
       tphhl$A1N$ZN = 1.0,
       tpllh$A2N$ZN = 1.0,
       tphhl$A2N$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tpllh$A1N$ZN$A2N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$A1N$ZN$A2N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tpllh$A1N$ZN$A2N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A1N$ZN$A2N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A1N$ZN$A2N_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A1N$ZN$A2N_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$A2N$ZN$A1N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$A2N$ZN$A1N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tpllh$A2N$ZN$A1N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A2N$ZN$A1N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A2N$ZN$A1N_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A2N$ZN$A1N_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1N_EQ_1_AN_A2N_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1N_EQ_1_AN_A2N_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$B2$ZN$A1N_EQ_1_AN_A2N_EQ_1_AN_B1_EQ_1 = 1.0,
       tphlh$B2$ZN$A1N_EQ_1_AN_A2N_EQ_1_AN_B1_EQ_1 = 1.0,
       tplhl$B2$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B1_EQ_1 = 1.0,
       tphlh$B2$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B1_EQ_1 = 1.0,
       tplhl$B2$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B1_EQ_1 = 1.0,
       tphlh$B2$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B1_EQ_1 = 1.0;

     // path delays
     if (A1N == 1'b1 && A2N == 1'b1 && B1 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1N_EQ_1_AN_A2N_EQ_1_AN_B1_EQ_1, tplhl$B2$ZN$A1N_EQ_1_AN_A2N_EQ_1_AN_B1_EQ_1);
     if (A1N == 1'b1 && A2N == 1'b0 && B1 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B1_EQ_1, tplhl$B2$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B1_EQ_1);
     if (A1N == 1'b0 && A2N == 1'b1 && B1 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B1_EQ_1, tplhl$B2$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B1_EQ_1);
     ifnone
       (B2 *> ZN) = (tphlh$B2$ZN,tplhl$B2$ZN);

     if (A1N == 1'b1 && A2N == 1'b1 && B2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1N_EQ_1_AN_A2N_EQ_1_AN_B2_EQ_1, tplhl$B1$ZN$A1N_EQ_1_AN_A2N_EQ_1_AN_B2_EQ_1);
     if (A1N == 1'b1 && A2N == 1'b0 && B2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B2_EQ_1, tplhl$B1$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B2_EQ_1);
     if (A1N == 1'b0 && A2N == 1'b1 && B2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B2_EQ_1, tplhl$B1$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B2_EQ_1);
     ifnone
       (B1 *> ZN) = (tphlh$B1$ZN,tplhl$B1$ZN);

     if (A1N == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A2N *> ZN) = (tpllh$A2N$ZN$A1N_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A2N$ZN$A1N_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1N == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A2N *> ZN) = (tpllh$A2N$ZN$A1N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A2N$ZN$A1N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A1N == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
       (A2N *> ZN) = (tpllh$A2N$ZN$A1N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0, tphhl$A2N$ZN$A1N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A2N *> ZN) = (tpllh$A2N$ZN,tphhl$A2N$ZN);

     if (A2N == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A1N *> ZN) = (tpllh$A1N$ZN$A2N_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A1N$ZN$A2N_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A2N == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A1N *> ZN) = (tpllh$A1N$ZN$A2N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A1N$ZN$A2N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A2N == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
       (A1N *> ZN) = (tpllh$A1N$ZN$A2N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0, tphhl$A1N$ZN$A2N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A1N *> ZN) = (tpllh$A1N$ZN,tphhl$A1N$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AON2BBD2 (ZN, A1N, A2N, B1, B2);
input  A1N ;
input  A2N ;
input  B1 ;
input  B2 ;
output ZN ;

   or  (I0_out, A1N, A2N);
   not (I1_out, I0_out);
   and (I2_out, B1, B2);
   or  (I3_out, I1_out, I2_out);
   not (ZN, I3_out);

   specify
     // delay parameters
     specparam
       tpllh$A1N$ZN = 1.0,
       tphhl$A1N$ZN = 1.0,
       tpllh$A2N$ZN = 1.0,
       tphhl$A2N$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tpllh$A1N$ZN$A2N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$A1N$ZN$A2N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tpllh$A1N$ZN$A2N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A1N$ZN$A2N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A1N$ZN$A2N_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A1N$ZN$A2N_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$A2N$ZN$A1N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$A2N$ZN$A1N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tpllh$A2N$ZN$A1N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A2N$ZN$A1N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A2N$ZN$A1N_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A2N$ZN$A1N_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1N_EQ_1_AN_A2N_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1N_EQ_1_AN_A2N_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$B2$ZN$A1N_EQ_1_AN_A2N_EQ_1_AN_B1_EQ_1 = 1.0,
       tphlh$B2$ZN$A1N_EQ_1_AN_A2N_EQ_1_AN_B1_EQ_1 = 1.0,
       tplhl$B2$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B1_EQ_1 = 1.0,
       tphlh$B2$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B1_EQ_1 = 1.0,
       tplhl$B2$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B1_EQ_1 = 1.0,
       tphlh$B2$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B1_EQ_1 = 1.0;

     // path delays
     if (A1N == 1'b1 && A2N == 1'b1 && B1 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1N_EQ_1_AN_A2N_EQ_1_AN_B1_EQ_1, tplhl$B2$ZN$A1N_EQ_1_AN_A2N_EQ_1_AN_B1_EQ_1);
     if (A1N == 1'b1 && A2N == 1'b0 && B1 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B1_EQ_1, tplhl$B2$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B1_EQ_1);
     if (A1N == 1'b0 && A2N == 1'b1 && B1 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B1_EQ_1, tplhl$B2$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B1_EQ_1);
     ifnone
       (B2 *> ZN) = (tphlh$B2$ZN,tplhl$B2$ZN);

     if (A1N == 1'b1 && A2N == 1'b1 && B2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1N_EQ_1_AN_A2N_EQ_1_AN_B2_EQ_1, tplhl$B1$ZN$A1N_EQ_1_AN_A2N_EQ_1_AN_B2_EQ_1);
     if (A1N == 1'b1 && A2N == 1'b0 && B2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B2_EQ_1, tplhl$B1$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B2_EQ_1);
     if (A1N == 1'b0 && A2N == 1'b1 && B2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B2_EQ_1, tplhl$B1$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B2_EQ_1);
     ifnone
       (B1 *> ZN) = (tphlh$B1$ZN,tplhl$B1$ZN);

     if (A1N == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A2N *> ZN) = (tpllh$A2N$ZN$A1N_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A2N$ZN$A1N_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1N == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A2N *> ZN) = (tpllh$A2N$ZN$A1N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A2N$ZN$A1N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A1N == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
       (A2N *> ZN) = (tpllh$A2N$ZN$A1N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0, tphhl$A2N$ZN$A1N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A2N *> ZN) = (tpllh$A2N$ZN,tphhl$A2N$ZN);

     if (A2N == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A1N *> ZN) = (tpllh$A1N$ZN$A2N_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A1N$ZN$A2N_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A2N == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A1N *> ZN) = (tpllh$A1N$ZN$A2N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A1N$ZN$A2N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A2N == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
       (A1N *> ZN) = (tpllh$A1N$ZN$A2N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0, tphhl$A1N$ZN$A2N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A1N *> ZN) = (tpllh$A1N$ZN,tphhl$A1N$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AON2BBD4 (ZN, A1N, A2N, B1, B2);
input  A1N ;
input  A2N ;
input  B1 ;
input  B2 ;
output ZN ;

   or  (I0_out, A1N, A2N);
   not (I1_out, I0_out);
   and (I2_out, B1, B2);
   or  (I3_out, I1_out, I2_out);
   not (ZN, I3_out);

   specify
     // delay parameters
     specparam
       tpllh$A1N$ZN = 1.0,
       tphhl$A1N$ZN = 1.0,
       tpllh$A2N$ZN = 1.0,
       tphhl$A2N$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tpllh$A1N$ZN$A2N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$A1N$ZN$A2N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tpllh$A1N$ZN$A2N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A1N$ZN$A2N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A1N$ZN$A2N_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A1N$ZN$A2N_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$A2N$ZN$A1N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$A2N$ZN$A1N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tpllh$A2N$ZN$A1N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A2N$ZN$A1N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A2N$ZN$A1N_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A2N$ZN$A1N_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1N_EQ_1_AN_A2N_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1N_EQ_1_AN_A2N_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$B2$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B1_EQ_1 = 1.0,
       tphlh$B2$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B1_EQ_1 = 1.0,
       tplhl$B2$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B1_EQ_1 = 1.0,
       tphlh$B2$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B1_EQ_1 = 1.0,
       tplhl$B2$ZN$A1N_EQ_1_AN_A2N_EQ_1_AN_B1_EQ_1 = 1.0,
       tphlh$B2$ZN$A1N_EQ_1_AN_A2N_EQ_1_AN_B1_EQ_1 = 1.0;

     // path delays
     if (A1N == 1'b1 && A2N == 1'b1 && B1 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1N_EQ_1_AN_A2N_EQ_1_AN_B1_EQ_1, tplhl$B2$ZN$A1N_EQ_1_AN_A2N_EQ_1_AN_B1_EQ_1);
     if (A1N == 1'b1 && A2N == 1'b0 && B1 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B1_EQ_1, tplhl$B2$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B1_EQ_1);
     if (A1N == 1'b0 && A2N == 1'b1 && B1 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B1_EQ_1, tplhl$B2$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B1_EQ_1);
     ifnone
       (B2 *> ZN) = (tphlh$B2$ZN,tplhl$B2$ZN);

     if (A1N == 1'b1 && A2N == 1'b1 && B2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1N_EQ_1_AN_A2N_EQ_1_AN_B2_EQ_1, tplhl$B1$ZN$A1N_EQ_1_AN_A2N_EQ_1_AN_B2_EQ_1);
     if (A1N == 1'b1 && A2N == 1'b0 && B2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B2_EQ_1, tplhl$B1$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B2_EQ_1);
     if (A1N == 1'b0 && A2N == 1'b1 && B2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B2_EQ_1, tplhl$B1$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B2_EQ_1);
     ifnone
       (B1 *> ZN) = (tphlh$B1$ZN,tplhl$B1$ZN);

     if (A1N == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A2N *> ZN) = (tpllh$A2N$ZN$A1N_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A2N$ZN$A1N_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1N == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A2N *> ZN) = (tpllh$A2N$ZN$A1N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A2N$ZN$A1N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A1N == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
       (A2N *> ZN) = (tpllh$A2N$ZN$A1N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0, tphhl$A2N$ZN$A1N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A2N *> ZN) = (tpllh$A2N$ZN,tphhl$A2N$ZN);

     if (A2N == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A1N *> ZN) = (tpllh$A1N$ZN$A2N_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A1N$ZN$A2N_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A2N == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A1N *> ZN) = (tpllh$A1N$ZN$A2N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A1N$ZN$A2N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A2N == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
       (A1N *> ZN) = (tpllh$A1N$ZN$A2N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0, tphhl$A1N$ZN$A2N_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A1N *> ZN) = (tpllh$A1N$ZN,tphhl$A1N$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AON2D1 (ZN, A1, A2, B1, B2);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
output ZN ;

   and (I0_out, B1, B2);
   and (I1_out, A1, A2);
   or  (I2_out, I0_out, I1_out);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1);
     ifnone
       (B2 *> ZN) = (tphlh$B2$ZN,tplhl$B2$ZN);

     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1);
     ifnone
       (B1 *> ZN) = (tphlh$B1$ZN,tplhl$B1$ZN);

     if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A2 *> ZN) = (tphlh$A2$ZN,tplhl$A2$ZN);

     if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A1 *> ZN) = (tphlh$A1$ZN,tplhl$A1$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AON2D2 (ZN, A1, A2, B1, B2);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
output ZN ;

   and (I0_out, A1, A2);
   and (I1_out, B1, B2);
   or  (I2_out, I0_out, I1_out);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1);
     ifnone
       (B2 *> ZN) = (tphlh$B2$ZN,tplhl$B2$ZN);

     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1);
     ifnone
       (B1 *> ZN) = (tphlh$B1$ZN,tplhl$B1$ZN);

     if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A2 *> ZN) = (tphlh$A2$ZN,tplhl$A2$ZN);

     if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A1 *> ZN) = (tphlh$A1$ZN,tplhl$A1$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AON2D4 (ZN, A1, A2, B1, B2);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
output ZN ;

   and (I0_out, A1, A2);
   and (I1_out, B1, B2);
   or  (I2_out, I0_out, I1_out);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1);
     ifnone
       (B2 *> ZN) = (tphlh$B2$ZN,tplhl$B2$ZN);

     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1);
     ifnone
       (B1 *> ZN) = (tphlh$B1$ZN,tplhl$B1$ZN);

     if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A2 *> ZN) = (tphlh$A2$ZN,tplhl$A2$ZN);

     if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A1 *> ZN) = (tphlh$A1$ZN,tplhl$A1$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AON3D1 (ZN, A1, A2, A3, B);
input  A1 ;
input  A2 ;
input  A3 ;
input  B ;
output ZN ;

   and (I1_out, A1, A2, A3);
   or  (I2_out, I1_out, B);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0,
       tplhl$B$ZN = 1.0,
       tphlh$B$ZN = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0 = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1 = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1 = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0);
     ifnone
       (B *> ZN) = (tphlh$B$ZN,tplhl$B$ZN);

     (A3 *> ZN) = (tphlh$A3$ZN, tplhl$A3$ZN);
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AON3D2 (ZN, A1, A2, A3, B);
input  A1 ;
input  A2 ;
input  A3 ;
input  B ;
output ZN ;

   and (I1_out, A1, A2, A3);
   or  (I2_out, I1_out, B);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0,
       tplhl$B$ZN = 1.0,
       tphlh$B$ZN = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0 = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1 = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1 = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0);
     ifnone
       (B *> ZN) = (tphlh$B$ZN,tplhl$B$ZN);

     (A3 *> ZN) = (tphlh$A3$ZN, tplhl$A3$ZN);
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AON3D4 (ZN, A1, A2, A3, B);
input  A1 ;
input  A2 ;
input  A3 ;
input  B ;
output ZN ;

   and (I1_out, A1, A2, A3);
   or  (I2_out, I1_out, B);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0,
       tplhl$B$ZN = 1.0,
       tphlh$B$ZN = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0 = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1 = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1 = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0);
     ifnone
       (B *> ZN) = (tphlh$B$ZN,tplhl$B$ZN);

     (A3 *> ZN) = (tphlh$A3$ZN, tplhl$A3$ZN);
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AON4D1 (ZN, A1, A2, A3, B1, B2);
input  A1 ;
input  A2 ;
input  A3 ;
input  B1 ;
input  B2 ;
output ZN ;

   and (I0_out, B1, B2);
   and (I2_out, A1, A2, A3);
   or  (I3_out, I0_out, I2_out);
   not (ZN, I3_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1);
     ifnone
       (B2 *> ZN) = (tphlh$B2$ZN,tplhl$B2$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_1, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_1, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_1, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_1, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_1);
     ifnone
       (B1 *> ZN) = (tphlh$B1$ZN,tplhl$B1$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A3 *> ZN) = (tphlh$A3$ZN,tplhl$A3$ZN);

     if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A2 *> ZN) = (tphlh$A2$ZN,tplhl$A2$ZN);

     if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A1 *> ZN) = (tphlh$A1$ZN,tplhl$A1$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AON4D2 (ZN, A1, A2, A3, B1, B2);
input  A1 ;
input  A2 ;
input  A3 ;
input  B1 ;
input  B2 ;
output ZN ;

   and (I1_out, A1, A2, A3);
   and (I2_out, B1, B2);
   or  (I3_out, I1_out, I2_out);
   not (ZN, I3_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1);
     ifnone
       (B2 *> ZN) = (tphlh$B2$ZN,tplhl$B2$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_1, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_1, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_1, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_1, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_1);
     ifnone
       (B1 *> ZN) = (tphlh$B1$ZN,tplhl$B1$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A3 *> ZN) = (tphlh$A3$ZN,tplhl$A3$ZN);

     if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A2 *> ZN) = (tphlh$A2$ZN,tplhl$A2$ZN);

     if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A1 *> ZN) = (tphlh$A1$ZN,tplhl$A1$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AON4D4 (ZN, A1, A2, A3, B1, B2);
input  A1 ;
input  A2 ;
input  A3 ;
input  B1 ;
input  B2 ;
output ZN ;

   and (I1_out, A1, A2, A3);
   and (I2_out, B1, B2);
   or  (I3_out, I1_out, I2_out);
   not (ZN, I3_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1);
     ifnone
       (B2 *> ZN) = (tphlh$B2$ZN,tplhl$B2$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_1, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_1, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_1, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_1, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_1);
     ifnone
       (B1 *> ZN) = (tphlh$B1$ZN,tplhl$B1$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A3 *> ZN) = (tphlh$A3$ZN,tplhl$A3$ZN);

     if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A2 *> ZN) = (tphlh$A2$ZN,tplhl$A2$ZN);

     if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A1 *> ZN) = (tphlh$A1$ZN,tplhl$A1$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AON5D1 (ZN, A1, A2, A3, B1, B2, B3);
input  A1 ;
input  A2 ;
input  A3 ;
input  B1 ;
input  B2 ;
input  B3 ;
output ZN ;

   and (I1_out, B1, B2, B3);
   and (I3_out, A1, A2, A3);
   or  (I4_out, I1_out, I3_out);
   not (ZN, I4_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tplhl$B3$ZN = 1.0,
       tphlh$B3$ZN = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$B3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$B3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$B3$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$B3$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$B3$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$B3$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$B3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$B3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (B3 *> ZN) = (tphlh$B3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tplhl$B3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
       (B3 *> ZN) = (tphlh$B3$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1, tplhl$B3$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
       (B3 *> ZN) = (tphlh$B3$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1, tplhl$B3$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (B3 *> ZN) = (tphlh$B3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tplhl$B3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     ifnone
       (B3 *> ZN) = (tphlh$B3$ZN,tplhl$B3$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1_AN_B3_EQ_1, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1_AN_B3_EQ_1, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B3_EQ_1, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B3_EQ_1, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B3_EQ_1);
     ifnone
       (B2 *> ZN) = (tphlh$B2$ZN,tplhl$B2$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1);
     ifnone
       (B1 *> ZN) = (tphlh$B1$ZN,tplhl$B1$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0, tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1, tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1, tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0, tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0);
     ifnone
       (A3 *> ZN) = (tphlh$A3$ZN,tplhl$A3$ZN);

     if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0);
     if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1, tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1);
     if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1, tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0);
     ifnone
       (A2 *> ZN) = (tphlh$A2$ZN,tplhl$A2$ZN);

     if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0);
     if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1, tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1);
     if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1, tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0);
     ifnone
       (A1 *> ZN) = (tphlh$A1$ZN,tplhl$A1$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AON5D2 (ZN, A1, A2, A3, B1, B2, B3);
input  A1 ;
input  A2 ;
input  A3 ;
input  B1 ;
input  B2 ;
input  B3 ;
output ZN ;

   and (I1_out, A1, A2, A3);
   and (I3_out, B1, B2, B3);
   or  (I4_out, I1_out, I3_out);
   not (ZN, I4_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tplhl$B3$ZN = 1.0,
       tphlh$B3$ZN = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$B3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$B3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$B3$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$B3$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$B3$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$B3$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$B3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$B3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (B3 *> ZN) = (tphlh$B3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tplhl$B3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
       (B3 *> ZN) = (tphlh$B3$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1, tplhl$B3$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
       (B3 *> ZN) = (tphlh$B3$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1, tplhl$B3$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (B3 *> ZN) = (tphlh$B3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tplhl$B3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     ifnone
       (B3 *> ZN) = (tphlh$B3$ZN,tplhl$B3$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1_AN_B3_EQ_1, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1_AN_B3_EQ_1, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B3_EQ_1, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B3_EQ_1, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B3_EQ_1);
     ifnone
       (B2 *> ZN) = (tphlh$B2$ZN,tplhl$B2$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1);
     ifnone
       (B1 *> ZN) = (tphlh$B1$ZN,tplhl$B1$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0, tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1, tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1, tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0, tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0);
     ifnone
       (A3 *> ZN) = (tphlh$A3$ZN,tplhl$A3$ZN);

     if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0);
     if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1, tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1);
     if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1, tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0);
     ifnone
       (A2 *> ZN) = (tphlh$A2$ZN,tplhl$A2$ZN);

     if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0);
     if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1, tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1);
     if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1, tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0);
     ifnone
       (A1 *> ZN) = (tphlh$A1$ZN,tplhl$A1$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AON5D4 (ZN, A1, A2, A3, B1, B2, B3);
input  A1 ;
input  A2 ;
input  A3 ;
input  B1 ;
input  B2 ;
input  B3 ;
output ZN ;

   and (I1_out, A1, A2, A3);
   and (I3_out, B1, B2, B3);
   or  (I4_out, I1_out, I3_out);
   not (ZN, I4_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tplhl$B3$ZN = 1.0,
       tphlh$B3$ZN = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$B3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$B3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$B3$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$B3$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$B3$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$B3$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$B3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$B3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (B3 *> ZN) = (tphlh$B3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tplhl$B3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
       (B3 *> ZN) = (tphlh$B3$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1, tplhl$B3$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
       (B3 *> ZN) = (tphlh$B3$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1, tplhl$B3$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (B3 *> ZN) = (tphlh$B3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tplhl$B3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     ifnone
       (B3 *> ZN) = (tphlh$B3$ZN,tplhl$B3$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1_AN_B3_EQ_1, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1_AN_B3_EQ_1, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B3_EQ_1, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B3_EQ_1, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B3_EQ_1);
     ifnone
       (B2 *> ZN) = (tphlh$B2$ZN,tplhl$B2$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1);
     ifnone
       (B1 *> ZN) = (tphlh$B1$ZN,tplhl$B1$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0, tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1, tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1, tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0, tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0);
     ifnone
       (A3 *> ZN) = (tphlh$A3$ZN,tplhl$A3$ZN);

     if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0);
     if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1, tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1);
     if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1, tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0);
     ifnone
       (A2 *> ZN) = (tphlh$A2$ZN,tplhl$A2$ZN);

     if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_0);
     if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1, tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_1);
     if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1, tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0);
     ifnone
       (A1 *> ZN) = (tphlh$A1$ZN,tplhl$A1$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AON6D1 (ZN, A1, A2, B, C);
input  A1 ;
input  A2 ;
input  B ;
input  C ;
output ZN ;

   and (I0_out, A1, A2);
   or  (I2_out, I0_out, B, C);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$B$ZN = 1.0,
       tphlh$B$ZN = 1.0,
       tplhl$C$ZN = 1.0,
       tphlh$C$ZN = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_C_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_C_EQ_0 = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_0 = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_0 = 1.0,
       tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_0 = 1.0,
       tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_0 = 1.0,
       tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B_EQ_0 = 1.0,
       tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B_EQ_0 = 1.0,
       tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B_EQ_0 = 1.0,
       tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b0)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B_EQ_0, tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b0)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B_EQ_0, tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b0)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_0, tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_0);
     ifnone
       (C *> ZN) = (tphlh$C$ZN,tplhl$C$ZN);

     if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_0, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_0, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && C == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_C_EQ_0, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_C_EQ_0);
     ifnone
       (B *> ZN) = (tphlh$B$ZN,tplhl$B$ZN);

     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AON6D2 (ZN, A1, A2, B, C);
input  A1 ;
input  A2 ;
input  B ;
input  C ;
output ZN ;

   and (I0_out, A1, A2);
   or  (I2_out, I0_out, B, C);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$B$ZN = 1.0,
       tphlh$B$ZN = 1.0,
       tplhl$C$ZN = 1.0,
       tphlh$C$ZN = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_C_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_C_EQ_0 = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_0 = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_0 = 1.0,
       tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_0 = 1.0,
       tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_0 = 1.0,
       tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B_EQ_0 = 1.0,
       tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B_EQ_0 = 1.0,
       tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B_EQ_0 = 1.0,
       tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b0)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B_EQ_0, tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b0)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B_EQ_0, tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b0)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_0, tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_0);
     ifnone
       (C *> ZN) = (tphlh$C$ZN,tplhl$C$ZN);

     if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_0, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_0, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && C == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_C_EQ_0, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_C_EQ_0);
     ifnone
       (B *> ZN) = (tphlh$B$ZN,tplhl$B$ZN);

     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AON6D4 (ZN, A1, A2, B, C);
input  A1 ;
input  A2 ;
input  B ;
input  C ;
output ZN ;

   and (I0_out, A1, A2);
   or  (I2_out, I0_out, B, C);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$B$ZN = 1.0,
       tphlh$B$ZN = 1.0,
       tplhl$C$ZN = 1.0,
       tphlh$C$ZN = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_C_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_C_EQ_0 = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_0 = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_0 = 1.0,
       tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_0 = 1.0,
       tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_0 = 1.0,
       tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B_EQ_0 = 1.0,
       tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B_EQ_0 = 1.0,
       tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B_EQ_0 = 1.0,
       tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b0)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B_EQ_0, tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b0)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B_EQ_0, tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b0)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_0, tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_0);
     ifnone
       (C *> ZN) = (tphlh$C$ZN,tplhl$C$ZN);

     if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_0, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_0, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && C == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_C_EQ_0, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_C_EQ_0);
     ifnone
       (B *> ZN) = (tphlh$B$ZN,tplhl$B$ZN);

     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AON7D1 (ZN, A1, A2, B1, B2, C);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
input  C ;
output ZN ;

   and (I0_out, A1, A2);
   and (I1_out, B1, B2);
   or  (I3_out, I0_out, I1_out, C);
   not (ZN, I3_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tplhl$C$ZN = 1.0,
       tphlh$C$ZN = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C_EQ_0 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_C_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_C_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C_EQ_0 = 1.0,
       tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0, tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (C *> ZN) = (tphlh$C$ZN,tplhl$C$ZN);

     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C_EQ_0, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C_EQ_0, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_C_EQ_0, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_C_EQ_0);
     ifnone
       (B2 *> ZN) = (tphlh$B2$ZN,tplhl$B2$ZN);

     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C_EQ_0, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C_EQ_0, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1_AN_C_EQ_0, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1_AN_C_EQ_0);
     ifnone
       (B1 *> ZN) = (tphlh$B1$ZN,tplhl$B1$ZN);

     if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_0);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_0);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C_EQ_0);
     ifnone
       (A2 *> ZN) = (tphlh$A2$ZN,tplhl$A2$ZN);

     if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_0);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_0);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C_EQ_0);
     ifnone
       (A1 *> ZN) = (tphlh$A1$ZN,tplhl$A1$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AON7D2 (ZN, A1, A2, B1, B2, C);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
input  C ;
output ZN ;

   and (I0_out, A1, A2);
   and (I1_out, B1, B2);
   or  (I3_out, I0_out, I1_out, C);
   not (ZN, I3_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tplhl$C$ZN = 1.0,
       tphlh$C$ZN = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C_EQ_0 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_C_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_C_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C_EQ_0 = 1.0,
       tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0, tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (C *> ZN) = (tphlh$C$ZN,tplhl$C$ZN);

     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C_EQ_0, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C_EQ_0, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_C_EQ_0, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_C_EQ_0);
     ifnone
       (B2 *> ZN) = (tphlh$B2$ZN,tplhl$B2$ZN);

     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C_EQ_0, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C_EQ_0, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1_AN_C_EQ_0, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1_AN_C_EQ_0);
     ifnone
       (B1 *> ZN) = (tphlh$B1$ZN,tplhl$B1$ZN);

     if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_0);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_0);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C_EQ_0);
     ifnone
       (A2 *> ZN) = (tphlh$A2$ZN,tplhl$A2$ZN);

     if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_0);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_0);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C_EQ_0);
     ifnone
       (A1 *> ZN) = (tphlh$A1$ZN,tplhl$A1$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AON7D4 (ZN, A1, A2, B1, B2, C);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
input  C ;
output ZN ;

   and (I0_out, A1, A2);
   and (I1_out, B1, B2);
   or  (I3_out, I0_out, I1_out, C);
   not (ZN, I3_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tplhl$C$ZN = 1.0,
       tphlh$C$ZN = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C_EQ_0 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_C_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_C_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C_EQ_0 = 1.0,
       tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0, tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (C *> ZN) = (tphlh$C$ZN,tplhl$C$ZN);

     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C_EQ_0, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C_EQ_0, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_C_EQ_0, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_C_EQ_0);
     ifnone
       (B2 *> ZN) = (tphlh$B2$ZN,tplhl$B2$ZN);

     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C_EQ_0, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C_EQ_0, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1_AN_C_EQ_0, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1_AN_C_EQ_0);
     ifnone
       (B1 *> ZN) = (tphlh$B1$ZN,tplhl$B1$ZN);

     if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_0);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_0);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C_EQ_0);
     ifnone
       (A2 *> ZN) = (tphlh$A2$ZN,tplhl$A2$ZN);

     if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_0);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_0);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C_EQ_0);
     ifnone
       (A1 *> ZN) = (tphlh$A1$ZN,tplhl$A1$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AON8D1 (ZN, A1, A2, B1, B2, C1, C2);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
input  C1 ;
input  C2 ;
output ZN ;

   and (I0_out, A1, A2);
   and (I1_out, C1, C2);
   and (I3_out, B1, B2);
   or  (I4_out, I0_out, I1_out, I3_out);
   not (ZN, I4_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tplhl$C1$ZN = 1.0,
       tphlh$C1$ZN = 1.0,
       tplhl$C2$ZN = 1.0,
       tphlh$C2$ZN = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_0 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$C1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$C1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_1 = 1.0,
       tphlh$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_1 = 1.0,
       tplhl$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_1 = 1.0,
       tphlh$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_1 = 1.0,
       tplhl$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$C2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_1 = 1.0,
       tphlh$C2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_1 = 1.0,
       tplhl$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1 = 1.0,
       tphlh$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1 = 1.0,
       tplhl$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1 = 1.0,
       tphlh$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1 = 1.0,
       tplhl$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1 = 1.0,
       tphlh$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1 = 1.0,
       tplhl$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1 = 1.0,
       tphlh$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
       (C2 *> ZN) = (tphlh$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1, tplhl$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
       (C2 *> ZN) = (tphlh$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1, tplhl$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
       (C2 *> ZN) = (tphlh$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1, tplhl$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
       (C2 *> ZN) = (tphlh$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1, tplhl$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
       (C2 *> ZN) = (tphlh$C2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_1, tplhl$C2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_1);
     ifnone
       (C2 *> ZN) = (tphlh$C2$ZN,tplhl$C2$ZN);

     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
       (C1 *> ZN) = (tphlh$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_1, tplhl$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
       (C1 *> ZN) = (tphlh$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_1, tplhl$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
       (C1 *> ZN) = (tphlh$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_1, tplhl$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
       (C1 *> ZN) = (tphlh$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_1, tplhl$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
       (C1 *> ZN) = (tphlh$C1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_C2_EQ_1, tplhl$C1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_C2_EQ_1);
     ifnone
       (C1 *> ZN) = (tphlh$C1$ZN,tplhl$C1$ZN);

     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_0, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_0);
     ifnone
       (B2 *> ZN) = (tphlh$B2$ZN,tplhl$B2$ZN);

     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_0, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_0);
     ifnone
       (B1 *> ZN) = (tphlh$B1$ZN,tplhl$B1$ZN);

     if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_0);
     ifnone
       (A2 *> ZN) = (tphlh$A2$ZN,tplhl$A2$ZN);

     if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_0);
     ifnone
       (A1 *> ZN) = (tphlh$A1$ZN,tplhl$A1$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AON8D2 (ZN, A1, A2, B1, B2, C1, C2);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
input  C1 ;
input  C2 ;
output ZN ;

   and (I0_out, C1, C2);
   and (I1_out, A1, A2);
   and (I3_out, B1, B2);
   or  (I4_out, I0_out, I1_out, I3_out);
   not (ZN, I4_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tplhl$C1$ZN = 1.0,
       tphlh$C1$ZN = 1.0,
       tplhl$C2$ZN = 1.0,
       tphlh$C2$ZN = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_0 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$C1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$C1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_1 = 1.0,
       tphlh$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_1 = 1.0,
       tplhl$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_1 = 1.0,
       tphlh$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_1 = 1.0,
       tplhl$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$C2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_1 = 1.0,
       tphlh$C2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_1 = 1.0,
       tplhl$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1 = 1.0,
       tphlh$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1 = 1.0,
       tplhl$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1 = 1.0,
       tphlh$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1 = 1.0,
       tplhl$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1 = 1.0,
       tphlh$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1 = 1.0,
       tplhl$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1 = 1.0,
       tphlh$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
       (C2 *> ZN) = (tphlh$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1, tplhl$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
       (C2 *> ZN) = (tphlh$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1, tplhl$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
       (C2 *> ZN) = (tphlh$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1, tplhl$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
       (C2 *> ZN) = (tphlh$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1, tplhl$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
       (C2 *> ZN) = (tphlh$C2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_1, tplhl$C2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_1);
     ifnone
       (C2 *> ZN) = (tphlh$C2$ZN,tplhl$C2$ZN);

     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
       (C1 *> ZN) = (tphlh$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_1, tplhl$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
       (C1 *> ZN) = (tphlh$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_1, tplhl$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
       (C1 *> ZN) = (tphlh$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_1, tplhl$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
       (C1 *> ZN) = (tphlh$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_1, tplhl$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
       (C1 *> ZN) = (tphlh$C1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_C2_EQ_1, tplhl$C1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_C2_EQ_1);
     ifnone
       (C1 *> ZN) = (tphlh$C1$ZN,tplhl$C1$ZN);

     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_0, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_0);
     ifnone
       (B2 *> ZN) = (tphlh$B2$ZN,tplhl$B2$ZN);

     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_0, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_0);
     ifnone
       (B1 *> ZN) = (tphlh$B1$ZN,tplhl$B1$ZN);

     if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_0);
     ifnone
       (A2 *> ZN) = (tphlh$A2$ZN,tplhl$A2$ZN);

     if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_0);
     ifnone
       (A1 *> ZN) = (tphlh$A1$ZN,tplhl$A1$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AON8D4 (ZN, A1, A2, B1, B2, C1, C2);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
input  C1 ;
input  C2 ;
output ZN ;

   and (I0_out, C1, C2);
   and (I1_out, A1, A2);
   and (I3_out, B1, B2);
   or  (I4_out, I0_out, I1_out, I3_out);
   not (ZN, I4_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tplhl$C1$ZN = 1.0,
       tphlh$C1$ZN = 1.0,
       tplhl$C2$ZN = 1.0,
       tphlh$C2$ZN = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_0 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$C1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$C1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_1 = 1.0,
       tphlh$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_1 = 1.0,
       tplhl$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_1 = 1.0,
       tphlh$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_1 = 1.0,
       tplhl$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$C2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_1 = 1.0,
       tphlh$C2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_1 = 1.0,
       tplhl$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1 = 1.0,
       tphlh$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1 = 1.0,
       tplhl$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1 = 1.0,
       tphlh$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1 = 1.0,
       tplhl$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1 = 1.0,
       tphlh$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1 = 1.0,
       tplhl$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1 = 1.0,
       tphlh$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
       (C2 *> ZN) = (tphlh$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1, tplhl$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
       (C2 *> ZN) = (tphlh$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1, tplhl$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
       (C2 *> ZN) = (tphlh$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1, tplhl$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
       (C2 *> ZN) = (tphlh$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1, tplhl$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
       (C2 *> ZN) = (tphlh$C2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_1, tplhl$C2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_1);
     ifnone
       (C2 *> ZN) = (tphlh$C2$ZN,tplhl$C2$ZN);

     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
       (C1 *> ZN) = (tphlh$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_1, tplhl$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
       (C1 *> ZN) = (tphlh$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_1, tplhl$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
       (C1 *> ZN) = (tphlh$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_1, tplhl$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
       (C1 *> ZN) = (tphlh$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_1, tplhl$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
       (C1 *> ZN) = (tphlh$C1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_C2_EQ_1, tplhl$C1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_C2_EQ_1);
     ifnone
       (C1 *> ZN) = (tphlh$C1$ZN,tplhl$C1$ZN);

     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_0, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_C1_EQ_0_AN_C2_EQ_0);
     ifnone
       (B2 *> ZN) = (tphlh$B2$ZN,tplhl$B2$ZN);

     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_0, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_0);
     ifnone
       (B1 *> ZN) = (tphlh$B1$ZN,tplhl$B1$ZN);

     if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_0);
     ifnone
       (A2 *> ZN) = (tphlh$A2$ZN,tplhl$A2$ZN);

     if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_0);
     ifnone
       (A1 *> ZN) = (tphlh$A1$ZN,tplhl$A1$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AX01D1 (Z, A1, A2, B);
input  A1 ;
input  A2 ;
input  B ;
output Z ;

   and (I0_out, A1, A2);
   xor (Z, I0_out, B);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tplhl$A1$Z = 1.0,
       tphlh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tplhl$A2$Z = 1.0,
       tphlh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$B$Z = 1.0,
       tplhl$B$Z = 1.0,
       tphlh$B$Z = 1.0,
       tphhl$B$Z = 1.0,
       tpllh$B$Z$A1_EQ_0_AN_A2_EQ_0 = 1.0,
       tphhl$B$Z$A1_EQ_0_AN_A2_EQ_0 = 1.0,
       tpllh$B$Z$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tphhl$B$Z$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tpllh$B$Z$A1_EQ_1_AN_A2_EQ_0 = 1.0,
       tphhl$B$Z$A1_EQ_1_AN_A2_EQ_0 = 1.0;

     // path delays
      (posedge B => (Z +: Z)) = (1.0, 1.0);
      (negedge B => (Z -: Z)) = (1.0, 1.0);

     if (A1 == 1'b1 && A2 == 1'b0)
       (B *> Z) = (tpllh$B$Z$A1_EQ_1_AN_A2_EQ_0, tphhl$B$Z$A1_EQ_1_AN_A2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1)
       (B *> Z) = (tpllh$B$Z$A1_EQ_0_AN_A2_EQ_1, tphhl$B$Z$A1_EQ_0_AN_A2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0)
       (B *> Z) = (tpllh$B$Z$A1_EQ_0_AN_A2_EQ_0, tphhl$B$Z$A1_EQ_0_AN_A2_EQ_0);
  //   ifnone
    //   (B *> Z) = (tpllh$B$Z,tplhl$B$Z);

     (posedge A2 *> (Z +: B^A1)) = (tpllh$A2$Z, tplhl$A2$Z);
     (negedge A2 *> (Z +: B)) = (tphlh$A2$Z, tphhl$A2$Z);
     (posedge A1 *> (Z +: B^A2)) = (tpllh$A1$Z, tplhl$A1$Z);
     (negedge A1 *> (Z +: B)) = (tphlh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AX01D2 (Z, A1, A2, B);
input  A1 ;
input  A2 ;
input  B ;
output Z ;

   and (I0_out, A1, A2);
   xor (Z, I0_out, B);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tplhl$A1$Z = 1.0,
       tphlh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tplhl$A2$Z = 1.0,
       tphlh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$B$Z = 1.0,
       tplhl$B$Z = 1.0,
       tphlh$B$Z = 1.0,
       tphhl$B$Z = 1.0,
       tpllh$B$Z$A1_EQ_0_AN_A2_EQ_0 = 1.0,
       tphhl$B$Z$A1_EQ_0_AN_A2_EQ_0 = 1.0,
       tpllh$B$Z$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tphhl$B$Z$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tpllh$B$Z$A1_EQ_1_AN_A2_EQ_0 = 1.0,
       tphhl$B$Z$A1_EQ_1_AN_A2_EQ_0 = 1.0;

   /*  // path delays
     if (A1 == 1'b1 && A2 == 1'b0)
       (B *> Z) = (tpllh$B$Z$A1_EQ_1_AN_A2_EQ_0, tphhl$B$Z$A1_EQ_1_AN_A2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1)
       (B *> Z) = (tpllh$B$Z$A1_EQ_0_AN_A2_EQ_1, tphhl$B$Z$A1_EQ_0_AN_A2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0)
       (B *> Z) = (tpllh$B$Z$A1_EQ_0_AN_A2_EQ_0, tphhl$B$Z$A1_EQ_0_AN_A2_EQ_0);
     ifnone
       (B *> Z) = (tpllh$B$Z,tplhl$B$Z);*/

     (posedge A2 *> (Z +: B^A1)) = (tpllh$A2$Z, tplhl$A2$Z);
     (negedge A2 *> (Z +: B)) = (tphlh$A2$Z, tphhl$A2$Z);
     (posedge A1 *> (Z +: B^A2)) = (tpllh$A1$Z, tplhl$A1$Z);
     (negedge A1 *> (Z +: B)) = (tphlh$A1$Z, tphhl$A1$Z);


      (posedge B => (Z +: Z)) = (1.0, 1.0);
      (negedge B => (Z -: Z)) = (1.0, 1.0);
      if (A1 == 1'b0 && A2 == 1'b0) (B +=> Z) = (1.0, 1.0);
      if (A1 == 1'b0 && A2 == 1'b1) (B +=> Z) = (1.0, 1.0);
      if (A1 == 1'b1 && A2 == 1'b0) (B +=> Z) = (1.0, 1.0);


   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AX01D4 (Z, A1, A2, B);
input  A1 ;
input  A2 ;
input  B ;
output Z ;

   and (I0_out, A1, A2);
   xor (Z, I0_out, B);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tplhl$A1$Z = 1.0,
       tphlh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tplhl$A2$Z = 1.0,
       tphlh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$B$Z = 1.0,
       tplhl$B$Z = 1.0,
       tphlh$B$Z = 1.0,
       tphhl$B$Z = 1.0,
       tpllh$B$Z$A1_EQ_0_AN_A2_EQ_0 = 1.0,
       tphhl$B$Z$A1_EQ_0_AN_A2_EQ_0 = 1.0,
       tpllh$B$Z$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tphhl$B$Z$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tpllh$B$Z$A1_EQ_1_AN_A2_EQ_0 = 1.0,
       tphhl$B$Z$A1_EQ_1_AN_A2_EQ_0 = 1.0;

     // path delays
 /*    if (A1 == 1'b1 && A2 == 1'b0)
       (B *> Z) = (tpllh$B$Z$A1_EQ_1_AN_A2_EQ_0, tphhl$B$Z$A1_EQ_1_AN_A2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1)
       (B *> Z) = (tpllh$B$Z$A1_EQ_0_AN_A2_EQ_1, tphhl$B$Z$A1_EQ_0_AN_A2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0)
       (B *> Z) = (tpllh$B$Z$A1_EQ_0_AN_A2_EQ_0, tphhl$B$Z$A1_EQ_0_AN_A2_EQ_0);
     ifnone
       (B *> Z) = (tpllh$B$Z,tplhl$B$Z);*/

     (posedge A2 *> (Z +: B^A1)) = (tpllh$A2$Z, tplhl$A2$Z);
     (negedge A2 *> (Z +: B)) = (tphlh$A2$Z, tphhl$A2$Z);
     (posedge A1 *> (Z +: B^A2)) = (tpllh$A1$Z, tplhl$A1$Z);
     (negedge A1 *> (Z +: B)) = (tphlh$A1$Z, tphhl$A1$Z);

      (posedge B => (Z +: Z)) = (1.0, 1.0);
      (negedge B => (Z -: Z)) = (1.0, 1.0);
      if (A1 == 1'b0 && A2 == 1'b0) (B +=> Z) = (1.0, 1.0);
      if (A1 == 1'b0 && A2 == 1'b1) (B +=> Z) = (1.0, 1.0);
      if (A1 == 1'b1 && A2 == 1'b0) (B +=> Z) = (1.0, 1.0);



   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AX02D1 (Z, A1, A2, B1, B2);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
output Z ;

   and (I0_out, B1, B2);
   and (I1_out, A1, A2);
   xor (Z, I0_out, I1_out);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tplhl$A1$Z = 1.0,
       tphlh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tplhl$A2$Z = 1.0,
       tphlh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$B1$Z = 1.0,
       tplhl$B1$Z = 1.0,
       tphlh$B1$Z = 1.0,
       tphhl$B1$Z = 1.0,
       tpllh$B2$Z = 1.0,
       tplhl$B2$Z = 1.0,
       tphlh$B2$Z = 1.0,
       tphhl$B2$Z = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1);
     ifnone
       (B2 *> Z) = (tpllh$B2$Z,tplhl$B2$Z);

     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1);
     ifnone
       (B1 *> Z) = (tpllh$B1$Z,tplhl$B1$Z);

     if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A2 *> Z) = (tpllh$A2$Z,tplhl$A2$Z);

     if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A1 *> Z) = (tpllh$A1$Z,tplhl$A1$Z);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AX02D2 (Z, A1, A2, B1, B2);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
output Z ;

   and (I0_out, B1, B2);
   and (I1_out, A1, A2);
   xor (Z, I0_out, I1_out);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tplhl$A1$Z = 1.0,
       tphlh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tplhl$A2$Z = 1.0,
       tphlh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$B1$Z = 1.0,
       tplhl$B1$Z = 1.0,
       tphlh$B1$Z = 1.0,
       tphhl$B1$Z = 1.0,
       tpllh$B2$Z = 1.0,
       tplhl$B2$Z = 1.0,
       tphlh$B2$Z = 1.0,
       tphhl$B2$Z = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1);
     ifnone
       (B2 *> Z) = (tpllh$B2$Z,tplhl$B2$Z);

     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1);
     ifnone
       (B1 *> Z) = (tpllh$B1$Z,tplhl$B1$Z);

     if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A2 *> Z) = (tpllh$A2$Z,tplhl$A2$Z);

     if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A1 *> Z) = (tpllh$A1$Z,tplhl$A1$Z);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AX02D4 (Z, A1, A2, B1, B2);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
output Z ;

   and (I0_out, B1, B2);
   and (I1_out, A1, A2);
   xor (Z, I0_out, I1_out);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tplhl$A1$Z = 1.0,
       tphlh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tplhl$A2$Z = 1.0,
       tphlh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$B1$Z = 1.0,
       tplhl$B1$Z = 1.0,
       tphlh$B1$Z = 1.0,
       tphhl$B1$Z = 1.0,
       tpllh$B2$Z = 1.0,
       tplhl$B2$Z = 1.0,
       tphlh$B2$Z = 1.0,
       tphhl$B2$Z = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1);
     ifnone
       (B2 *> Z) = (tpllh$B2$Z,tplhl$B2$Z);

     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1);
     ifnone
       (B1 *> Z) = (tpllh$B1$Z,tplhl$B1$Z);

     if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tphhl$A2$Z$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A2 *> Z) = (tpllh$A2$Z,tplhl$A2$Z);

     if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tphhl$A1$Z$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A1 *> Z) = (tpllh$A1$Z,tplhl$A1$Z);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AXN1D1 (ZN, A1, A2, B);
input  A1 ;
input  A2 ;
input  B ;
output ZN ;

   and (I0_out, A1, A2);
   xor (I1_out, I0_out, B);
   not (ZN, I1_out);

   specify
     // delay parameters
     specparam
       tpllh$A1$ZN = 1.0,
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tphhl$A1$ZN = 1.0,
       tpllh$A2$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tphhl$A2$ZN = 1.0,
       tpllh$B$ZN = 1.0,
       tplhl$B$ZN = 1.0,
       tphlh$B$ZN = 1.0,
       tphhl$B$ZN = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_0 = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0;

     // path delays
 /*    if (A1 == 1'b1 && A2 == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_0, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_0);
     ifnone
       (B *> ZN) = (tpllh$B$ZN,tplhl$B$ZN);*/

      (posedge B => (ZN +: ZN)) = (1.0, 1.0);
      (negedge B => (ZN -: ZN)) = (1.0, 1.0);
      if (A1 == 1'b0 && A2 == 1'b0) (B -=> ZN) = (1.0, 1.0);
      if (A1 == 1'b1 && A2 == 1'b0) (B -=> ZN) = (1.0, 1.0);
      if (A1 == 1'b0 && A2 == 1'b1) (B -=> ZN) = (1.0, 1.0);


     (posedge A2 *> (ZN +: !(B^A1))) = (tpllh$A2$ZN, tplhl$A2$ZN);
     (negedge A2 *> (ZN +: !B)) = (tphlh$A2$ZN, tphhl$A2$ZN);
     (posedge A1 *> (ZN +: !(B^A2))) = (tpllh$A1$ZN, tplhl$A1$ZN);
     (negedge A1 *> (ZN +: !B)) = (tphlh$A1$ZN, tphhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AXN1D2 (ZN, A1, A2, B);
input  A1 ;
input  A2 ;
input  B ;
output ZN ;

   and (I0_out, A1, A2);
   xor (I1_out, I0_out, B);
   not (ZN, I1_out);

   specify
     // delay parameters
     specparam
       tpllh$A1$ZN = 1.0,
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tphhl$A1$ZN = 1.0,
       tpllh$A2$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tphhl$A2$ZN = 1.0,
       tpllh$B$ZN = 1.0,
       tplhl$B$ZN = 1.0,
       tphlh$B$ZN = 1.0,
       tphhl$B$ZN = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_0 = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0;

     // path delays
/*     if (A1 == 1'b1 && A2 == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_0, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_0);
     ifnone
       (B *> ZN) = (tpllh$B$ZN,tplhl$B$ZN);*/


      (posedge B => (ZN +: ZN)) = (1.0, 1.0);
      (negedge B => (ZN -: ZN)) = (1.0, 1.0);
      if (A1 == 1'b0 && A2 == 1'b0) (B -=> ZN) = (1.0, 1.0);
      if (A1 == 1'b1 && A2 == 1'b0) (B -=> ZN) = (1.0, 1.0);
      if (A1 == 1'b0 && A2 == 1'b1) (B -=> ZN) = (1.0, 1.0);


     (posedge A2 *> (ZN +: !(B^A1))) = (tpllh$A2$ZN, tplhl$A2$ZN);
     (negedge A2 *> (ZN +: !B)) = (tphlh$A2$ZN, tphhl$A2$ZN);
     (posedge A1 *> (ZN +: !(B^A2))) = (tpllh$A1$ZN, tplhl$A1$ZN);
     (negedge A1 *> (ZN +: !B)) = (tphlh$A1$ZN, tphhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AXN1D4 (ZN, A1, A2, B);
input  A1 ;
input  A2 ;
input  B ;
output ZN ;

   and (I0_out, A1, A2);
   xor (I1_out, I0_out, B);
   not (ZN, I1_out);

   specify
     // delay parameters
     specparam
       tpllh$A1$ZN = 1.0,
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tphhl$A1$ZN = 1.0,
       tpllh$A2$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tphhl$A2$ZN = 1.0,
       tpllh$B$ZN = 1.0,
       tplhl$B$ZN = 1.0,
       tphlh$B$ZN = 1.0,
       tphhl$B$ZN = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_0 = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0;

     // path delays
 /*    if (A1 == 1'b1 && A2 == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_0, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_0);
     ifnone
       (B *> ZN) = (tpllh$B$ZN,tplhl$B$ZN);*/


      (posedge B => (ZN +: ZN)) = (1.0, 1.0);
      (negedge B => (ZN -: ZN)) = (1.0, 1.0);
      if (A1 == 1'b0 && A2 == 1'b0) (B -=> ZN) = (1.0, 1.0);
      if (A1 == 1'b1 && A2 == 1'b0) (B -=> ZN) = (1.0, 1.0);
      if (A1 == 1'b0 && A2 == 1'b1) (B -=> ZN) = (1.0, 1.0);

     (posedge A2 *> (ZN +: !(B^A1))) = (tpllh$A2$ZN, tplhl$A2$ZN);
     (negedge A2 *> (ZN +: !B)) = (tphlh$A2$ZN, tphhl$A2$ZN);
     (posedge A1 *> (ZN +: !(B^A2))) = (tpllh$A1$ZN, tplhl$A1$ZN);
     (negedge A1 *> (ZN +: !B)) = (tphlh$A1$ZN, tphhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AXN2D1 (ZN, A1, A2, B1, B2);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
output ZN ;

   and (I0_out, A1, A2);
   and (I1_out, B1, B2);
   xor (I2_out, I0_out, I1_out);
   not (ZN, I2_out);

   specify
     // delay parameters
 /*    specparam
       tpllh$A1$ZN = 1.0,
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tphhl$A1$ZN = 1.0,
       tpllh$A2$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tphhl$A2$ZN = 1.0,
       tpllh$B1$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tphhl$B1$ZN = 1.0,
       tpllh$B2$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tphhl$B2$ZN = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1);
     ifnone
       (B2 *> ZN) = (tpllh$B2$ZN,tplhl$B2$ZN);

     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1);
     ifnone
       (B1 *> ZN) = (tpllh$B1$ZN,tplhl$B1$ZN);

     if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A2 *> ZN) = (tpllh$A2$ZN,tplhl$A2$ZN);

     if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A1 *> ZN) = (tpllh$A1$ZN,tplhl$A1$ZN);*/

      (posedge A1 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge A1 => (ZN -: ZN)) = (1.0, 1.0);
      if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0) (A1 -=> ZN) = (1.0, 1.0);
      if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1) (A1 -=> ZN) = (1.0, 1.0);
      if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0) (A1 -=> ZN) = (1.0, 1.0);
     
      (posedge A2 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge A2 => (ZN -: ZN)) = (1.0, 1.0);
      if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0) (A2 -=> ZN) = (1.0, 1.0);
      if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0) (A2 -=> ZN) = (1.0, 1.0);
      if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1) (A2 -=> ZN) = (1.0, 1.0);

      (posedge B1 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge B1 => (ZN -: ZN)) = (1.0, 1.0);
      if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1) (B1 -=> ZN) = (1.0, 1.0);
      if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1) (B1 -=> ZN) = (1.0, 1.0);
      if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1) (B1 -=> ZN) = (1.0, 1.0);
     
     
      (posedge B2 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge B2 => (ZN -: ZN)) = (1.0, 1.0);
      if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1) (B2 -=> ZN) = (1.0, 1.0);
      if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1) (B2 -=> ZN) = (1.0, 1.0);
      if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1) (B2 -=> ZN) = (1.0, 1.0);


   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AXN2D2 (ZN, A1, A2, B1, B2);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
output ZN ;

   and (I0_out, A1, A2);
   and (I1_out, B1, B2);
   xor (I2_out, I0_out, I1_out);
   not (ZN, I2_out);

   specify
     // delay parameters
/*     specparam
       tpllh$A1$ZN = 1.0,
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tphhl$A1$ZN = 1.0,
       tpllh$A2$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tphhl$A2$ZN = 1.0,
       tpllh$B1$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tphhl$B1$ZN = 1.0,
       tpllh$B2$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tphhl$B2$ZN = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1);
     ifnone
       (B2 *> ZN) = (tpllh$B2$ZN,tplhl$B2$ZN);

     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1);
     ifnone
       (B1 *> ZN) = (tpllh$B1$ZN,tplhl$B1$ZN);

     if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A2 *> ZN) = (tpllh$A2$ZN,tplhl$A2$ZN);

     if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A1 *> ZN) = (tpllh$A1$ZN,tplhl$A1$ZN);*/


      (posedge A1 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge A1 => (ZN -: ZN)) = (1.0, 1.0);
      if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0) (A1 -=> ZN) = (1.0, 1.0);
      if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1) (A1 -=> ZN) = (1.0, 1.0);
      if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0) (A1 -=> ZN) = (1.0, 1.0);
     
      (posedge A2 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge A2 => (ZN -: ZN)) = (1.0, 1.0);
      if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0) (A2 -=> ZN) = (1.0, 1.0);
      if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0) (A2 -=> ZN) = (1.0, 1.0);
      if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1) (A2 -=> ZN) = (1.0, 1.0);

      (posedge B1 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge B1 => (ZN -: ZN)) = (1.0, 1.0);
      if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1) (B1 -=> ZN) = (1.0, 1.0);
      if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1) (B1 -=> ZN) = (1.0, 1.0);
      if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1) (B1 -=> ZN) = (1.0, 1.0);
     
     
      (posedge B2 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge B2 => (ZN -: ZN)) = (1.0, 1.0);
      if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1) (B2 -=> ZN) = (1.0, 1.0);
      if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1) (B2 -=> ZN) = (1.0, 1.0);
      if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1) (B2 -=> ZN) = (1.0, 1.0);


   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_AXN2D4 (ZN, A1, A2, B1, B2);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
output ZN ;

   and (I0_out, A1, A2);
   and (I1_out, B1, B2);
   xor (I2_out, I0_out, I1_out);
   not (ZN, I2_out);

   specify
     // delay parameters
/*     specparam
       tpllh$A1$ZN = 1.0,
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tphhl$A1$ZN = 1.0,
       tpllh$A2$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tphhl$A2$ZN = 1.0,
       tpllh$B1$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tphhl$B1$ZN = 1.0,
       tpllh$B2$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tphhl$B2$ZN = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1);
     ifnone
       (B2 *> ZN) = (tpllh$B2$ZN,tplhl$B2$ZN);

     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B2_EQ_1);
     ifnone
       (B1 *> ZN) = (tpllh$B1$ZN,tplhl$B1$ZN);

     if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tplhl$A2$ZN$A1_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A2 *> ZN) = (tpllh$A2$ZN,tplhl$A2$ZN);

     if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tplhl$A1$ZN$A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (A1 *> ZN) = (tpllh$A1$ZN,tplhl$A1$ZN);*/

      (posedge A1 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge A1 => (ZN -: ZN)) = (1.0, 1.0);
      if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0) (A1 -=> ZN) = (1.0, 1.0);
      if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1) (A1 -=> ZN) = (1.0, 1.0);
      if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0) (A1 -=> ZN) = (1.0, 1.0);
     
      (posedge A2 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge A2 => (ZN -: ZN)) = (1.0, 1.0);
      if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0) (A2 -=> ZN) = (1.0, 1.0);
      if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0) (A2 -=> ZN) = (1.0, 1.0);
      if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1) (A2 -=> ZN) = (1.0, 1.0);

      (posedge B1 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge B1 => (ZN -: ZN)) = (1.0, 1.0);
      if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1) (B1 -=> ZN) = (1.0, 1.0);
      if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1) (B1 -=> ZN) = (1.0, 1.0);
      if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1) (B1 -=> ZN) = (1.0, 1.0);
     
     
      (posedge B2 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge B2 => (ZN -: ZN)) = (1.0, 1.0);
      if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1) (B2 -=> ZN) = (1.0, 1.0);
      if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1) (B2 -=> ZN) = (1.0, 1.0);
      if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1) (B2 -=> ZN) = (1.0, 1.0);





   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_BF01D1 (Z, I);
input  I ;
output Z ;

   buf (Z, I);

   specify
     // delay parameters
     specparam
       tpllh$I$Z = 1.0,
       tphhl$I$Z = 1.0;

     // path delays
     (I *> Z) = (tpllh$I$Z, tphhl$I$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_BF01D12 (Z, I);
input  I ;
output Z ;

   buf (Z, I);

   specify
     // delay parameters
     specparam
       tpllh$I$Z = 1.0,
       tphhl$I$Z = 1.0;

     // path delays
     (I *> Z) = (tpllh$I$Z, tphhl$I$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_BF01D16 (Z, I);
input  I ;
output Z ;

   buf (Z, I);

   specify
     // delay parameters
     specparam
       tpllh$I$Z = 1.0,
       tphhl$I$Z = 1.0;

     // path delays
     (I *> Z) = (tpllh$I$Z, tphhl$I$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_BF01D2 (Z, I);
input  I ;
output Z ;

   buf (Z, I);

   specify
     // delay parameters
     specparam
       tpllh$I$Z = 1.0,
       tphhl$I$Z = 1.0;

     // path delays
     (I *> Z) = (tpllh$I$Z, tphhl$I$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_BF01D20 (Z, I);
input  I ;
output Z ;

   buf (Z, I);

   specify
     // delay parameters
     specparam
       tpllh$I$Z = 1.0,
       tphhl$I$Z = 1.0;

     // path delays
     (I *> Z) = (tpllh$I$Z, tphhl$I$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_BF01D3 (Z, I);
input  I ;
output Z ;

   buf (Z, I);

   specify
     // delay parameters
     specparam
       tpllh$I$Z = 1.0,
       tphhl$I$Z = 1.0;

     // path delays
     (I *> Z) = (tpllh$I$Z, tphhl$I$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_BF01D4 (Z, I);
input  I ;
output Z ;

   buf (Z, I);

   specify
     // delay parameters
     specparam
       tpllh$I$Z = 1.0,
       tphhl$I$Z = 1.0;

     // path delays
     (I *> Z) = (tpllh$I$Z, tphhl$I$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_BF01D6 (Z, I);
input  I ;
output Z ;

   buf (Z, I);

   specify
     // delay parameters
     specparam
       tpllh$I$Z = 1.0,
       tphhl$I$Z = 1.0;

     // path delays
     (I *> Z) = (tpllh$I$Z, tphhl$I$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_BF01D8 (Z, I);
input  I ;
output Z ;

   buf (Z, I);

   specify
     // delay parameters
     specparam
       tpllh$I$Z = 1.0,
       tphhl$I$Z = 1.0;

     // path delays
     (I *> Z) = (tpllh$I$Z, tphhl$I$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_BH01D0 (D);
inout  D ;

   buf (weak1, weak0) (D, D);


endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
//`ifdef RST
module RT8_DF01D1 (Q, QN, CP, D);
input  CP ;
input  D ;
output Q ;
output QN ;
reg NOTIFIER ;
    reg ReSeT;
`ifdef  RSTn_lib

	 initial begin
		ReSeT = 0 ;
		#3 ReSeT = 1 ;
		#111 ReSeT = 0 ;
	end

  `else initial  ReSeT = 0;
//udp_dff (N_S_XM19_G, D, CP, 1'B0, 1'B0, NOTIFIER);
`endif



   udp_dff (N_S_XM19_G, D, CP, ReSeT /*1'B0*/, 1'B0, NOTIFIER);
   not (N_NET0130_XM16_D, N_S_XM19_G);
   buf (Q, N_S_XM19_G);
   not (QN, N_S_XM19_G);

   specify
     // delay parameters
     specparam
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tpllh$CP$QN = 1.0,
       tplhl$CP$QN = 1.0,
       tminpwh$CP$D_EQ_0 = 1.0,
       tminpwl$CP$D_EQ_0 = 1.0,
       tsetup_negedge$D$CP = 1.0,
       thold_negedge$D$CP = 1.0,
       tsetup_posedge$D$CP = 1.0,
       thold_posedge$D$CP = 1.0;

     // path delays
     (posedge CP *> (QN -: D)) = (tpllh$CP$QN, tplhl$CP$QN);
     (posedge CP *> (Q +: D)) = (tpllh$CP$Q, tplhl$CP$Q);
     $setuphold(posedge CP, negedge D, tsetup_negedge$D$CP, thold_negedge$D$CP, NOTIFIER);
     $setuphold(posedge CP, posedge D, tsetup_posedge$D$CP, thold_posedge$D$CP, NOTIFIER);
     $width(posedge CP &&& D == 1'b0, tminpwh$CP$D_EQ_0, 0, NOTIFIER);
     $width(negedge CP &&& D == 1'b0, tminpwl$CP$D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF01D2 (Q, QN, CP, D);
input  CP ;
input  D ;
output Q ;
output QN ;
reg NOTIFIER ;
reg ReSeT;

`ifdef  RSTn_lib

	 initial begin
		ReSeT = 0 ;
		#3 ReSeT = 1 ;
		#111 ReSeT = 0 ;
	end

  `else initial  ReSeT = 0;
//udp_dff (N_S_XM19_G, D, CP, 1'B0, 1'B0, NOTIFIER);
`endif



   udp_dff (N_S_XM19_G, D, CP, ReSeT, 1'B0, NOTIFIER);
   not (N_NET0130_XM16_D, N_S_XM19_G);
   buf (Q, N_S_XM19_G);
   not (QN, N_S_XM19_G);

   specify
     // delay parameters
     specparam
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tpllh$CP$QN = 1.0,
       tplhl$CP$QN = 1.0,
       tminpwh$CP$D_EQ_0 = 1.0,
       tminpwl$CP$D_EQ_0 = 1.0,
       tsetup_negedge$D$CP = 1.0,
       thold_negedge$D$CP = 1.0,
       tsetup_posedge$D$CP = 1.0,
       thold_posedge$D$CP = 1.0;

     // path delays
     (posedge CP *> (QN -: D)) = (tpllh$CP$QN, tplhl$CP$QN);
     (posedge CP *> (Q +: D)) = (tpllh$CP$Q, tplhl$CP$Q);
     $setuphold(posedge CP, negedge D, tsetup_negedge$D$CP, thold_negedge$D$CP, NOTIFIER);
     $setuphold(posedge CP, posedge D, tsetup_posedge$D$CP, thold_posedge$D$CP, NOTIFIER);
     $width(posedge CP &&& D == 1'b0, tminpwh$CP$D_EQ_0, 0, NOTIFIER);
     $width(negedge CP &&& D == 1'b0, tminpwl$CP$D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF01D4 (Q, QN, CP, D);
input  CP ;
input  D ;
output Q ;
output QN ;
reg NOTIFIER ;
reg ReSeT;

`ifdef  RSTn_lib
	 initial begin
		ReSeT = 0 ;
		#3 ReSeT = 1 ;
		#111 ReSeT = 0 ;
	end

  `else initial  ReSeT = 0;
`endif
udp_dff (N_S_XM19_G, D, CP, ReSeT /*1'B0*/, 1'B0, NOTIFIER);
   not (N_NET0130_XM16_D, N_S_XM19_G);
   buf (Q, N_S_XM19_G);
   not (QN, N_S_XM19_G);

   specify
     // delay parameters
     specparam
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tpllh$CP$QN = 1.0,
       tplhl$CP$QN = 1.0,
       tminpwh$CP$D_EQ_0 = 1.0,
       tminpwl$CP$D_EQ_0 = 1.0,
       tsetup_negedge$D$CP = 1.0,
       thold_negedge$D$CP = 1.0,
       tsetup_posedge$D$CP = 1.0,
       thold_posedge$D$CP = 1.0;

     // path delays
     (posedge CP *> (QN -: D)) = (tpllh$CP$QN, tplhl$CP$QN);
     (posedge CP *> (Q +: D)) = (tpllh$CP$Q, tplhl$CP$Q);
     $setuphold(posedge CP, negedge D, tsetup_negedge$D$CP, thold_negedge$D$CP, NOTIFIER);
     $setuphold(posedge CP, posedge D, tsetup_posedge$D$CP, thold_posedge$D$CP, NOTIFIER);
     $width(posedge CP &&& D == 1'b0, tminpwh$CP$D_EQ_0, 0, NOTIFIER);
     $width(negedge CP &&& D == 1'b0, tminpwl$CP$D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF01ED1 (Q, QN, CP, D, E);
input  CP ;
input  D ;
input  E ;
output Q ;
output QN ;
reg NOTIFIER ;

   udp_mux2 (I0_D, N_S_XM3_G, D, E);
   udp_dff (N_S_XM3_G, I0_D, CP, 1'B0, 1'B0, NOTIFIER);
   not (N_NET0235_XM29_G, N_S_XM3_G);
   not (Q, N_NET0235_XM29_G);
   buf (QN, N_NET0235_XM29_G);
   not (I7_out, D);
   and (D_EQ_0_AN_E_EQ_1, I7_out, E);

   specify
     // delay parameters
     specparam
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tpllh$CP$QN = 1.0,
       tplhl$CP$QN = 1.0,
       tminpwh$CP$D_EQ_0_AN_E_EQ_1 = 1.0,
       tminpwl$CP$D_EQ_0_AN_E_EQ_1 = 1.0,
       tsetup_negedge$D$CP$E_EQ_1 = 1.0,
       thold_negedge$D$CP$E_EQ_1 = 1.0,
       tsetup_negedge$E$CP$D_EQ_0 = 1.0,
       thold_negedge$E$CP$D_EQ_0 = 1.0,
       tsetup_negedge$E$CP$D_EQ_1 = 1.0,
       thold_negedge$E$CP$D_EQ_1 = 1.0,
       tsetup_posedge$D$CP$E_EQ_1 = 1.0,
       thold_posedge$D$CP$E_EQ_1 = 1.0,
       tsetup_posedge$E$CP$D_EQ_0 = 1.0,
       thold_posedge$E$CP$D_EQ_0 = 1.0,
       tsetup_posedge$E$CP$D_EQ_1 = 1.0,
       thold_posedge$E$CP$D_EQ_1 = 1.0;

     // path delays
     (posedge CP *> (QN -: E?D:N_S_XM3_G)) = (tpllh$CP$QN, tplhl$CP$QN);
     (posedge CP *> (Q +: E?D:N_S_XM3_G)) = (tpllh$CP$Q, tplhl$CP$Q);
     $setuphold(posedge CP &&& E == 1'b1, negedge D, tsetup_negedge$D$CP$E_EQ_1, thold_negedge$D$CP$E_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& D == 1'b0, negedge E, tsetup_negedge$E$CP$D_EQ_0, thold_negedge$E$CP$D_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& D == 1'b1, negedge E, tsetup_negedge$E$CP$D_EQ_1, thold_negedge$E$CP$D_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& E == 1'b1, posedge D, tsetup_posedge$D$CP$E_EQ_1, thold_posedge$D$CP$E_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& D == 1'b0, posedge E, tsetup_posedge$E$CP$D_EQ_0, thold_posedge$E$CP$D_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& D == 1'b1, posedge E, tsetup_posedge$E$CP$D_EQ_1, thold_posedge$E$CP$D_EQ_1, NOTIFIER);
     $width(posedge CP &&& D_EQ_0_AN_E_EQ_1 == 1'b1, tminpwh$CP$D_EQ_0_AN_E_EQ_1, 0, NOTIFIER);
     $width(negedge CP &&& D_EQ_0_AN_E_EQ_1 == 1'b1, tminpwl$CP$D_EQ_0_AN_E_EQ_1, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF01ED2 (Q, QN, CP, D, E);
input  CP ;
input  D ;
input  E ;
output Q ;
output QN ;
reg NOTIFIER ;

   udp_mux2 (I0_D, N_S_XM3_G, D, E);
   udp_dff (N_S_XM3_G, I0_D, CP, 1'B0, 1'B0, NOTIFIER);
   not (N_NET0235_XM29_G, N_S_XM3_G);
   not (Q, N_NET0235_XM29_G);
   buf (QN, N_NET0235_XM29_G);
   not (I7_out, D);
   and (D_EQ_0_AN_E_EQ_1, I7_out, E);

   specify
     // delay parameters
     specparam
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tpllh$CP$QN = 1.0,
       tplhl$CP$QN = 1.0,
       tminpwh$CP$D_EQ_0_AN_E_EQ_1 = 1.0,
       tminpwl$CP$D_EQ_0_AN_E_EQ_1 = 1.0,
       tsetup_negedge$D$CP$E_EQ_1 = 1.0,
       thold_negedge$D$CP$E_EQ_1 = 1.0,
       tsetup_negedge$E$CP$D_EQ_0 = 1.0,
       thold_negedge$E$CP$D_EQ_0 = 1.0,
       tsetup_negedge$E$CP$D_EQ_1 = 1.0,
       thold_negedge$E$CP$D_EQ_1 = 1.0,
       tsetup_posedge$D$CP$E_EQ_1 = 1.0,
       thold_posedge$D$CP$E_EQ_1 = 1.0,
       tsetup_posedge$E$CP$D_EQ_0 = 1.0,
       thold_posedge$E$CP$D_EQ_0 = 1.0,
       tsetup_posedge$E$CP$D_EQ_1 = 1.0,
       thold_posedge$E$CP$D_EQ_1 = 1.0;

     // path delays
     (posedge CP *> (QN -: E?D:N_S_XM3_G)) = (tpllh$CP$QN, tplhl$CP$QN);
     (posedge CP *> (Q +: E?D:N_S_XM3_G)) = (tpllh$CP$Q, tplhl$CP$Q);
     $setuphold(posedge CP &&& E == 1'b1, negedge D, tsetup_negedge$D$CP$E_EQ_1, thold_negedge$D$CP$E_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& D == 1'b0, negedge E, tsetup_negedge$E$CP$D_EQ_0, thold_negedge$E$CP$D_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& D == 1'b1, negedge E, tsetup_negedge$E$CP$D_EQ_1, thold_negedge$E$CP$D_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& E == 1'b1, posedge D, tsetup_posedge$D$CP$E_EQ_1, thold_posedge$D$CP$E_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& D == 1'b0, posedge E, tsetup_posedge$E$CP$D_EQ_0, thold_posedge$E$CP$D_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& D == 1'b1, posedge E, tsetup_posedge$E$CP$D_EQ_1, thold_posedge$E$CP$D_EQ_1, NOTIFIER);
     $width(posedge CP &&& D_EQ_0_AN_E_EQ_1 == 1'b1, tminpwh$CP$D_EQ_0_AN_E_EQ_1, 0, NOTIFIER);
     $width(negedge CP &&& D_EQ_0_AN_E_EQ_1 == 1'b1, tminpwl$CP$D_EQ_0_AN_E_EQ_1, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF01ED4 (Q, QN, CP, D, E);
input  CP ;
input  D ;
input  E ;
output Q ;
output QN ;
reg NOTIFIER ;

   udp_mux2 (I0_D, N_S_XM3_G, D, E);
   udp_dff (N_S_XM3_G, I0_D, CP, 1'B0, 1'B0, NOTIFIER);
   not (N_NET0235_XM29_G, N_S_XM3_G);
   not (Q, N_NET0235_XM29_G);
   buf (QN, N_NET0235_XM29_G);
   not (I7_out, D);
   and (D_EQ_0_AN_E_EQ_1, I7_out, E);

   specify
     // delay parameters
     specparam
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tpllh$CP$QN = 1.0,
       tplhl$CP$QN = 1.0,
       tminpwh$CP$D_EQ_0_AN_E_EQ_1 = 1.0,
       tminpwl$CP$D_EQ_0_AN_E_EQ_1 = 1.0,
       tsetup_negedge$D$CP$E_EQ_1 = 1.0,
       thold_negedge$D$CP$E_EQ_1 = 1.0,
       tsetup_negedge$E$CP$D_EQ_0 = 1.0,
       thold_negedge$E$CP$D_EQ_0 = 1.0,
       tsetup_negedge$E$CP$D_EQ_1 = 1.0,
       thold_negedge$E$CP$D_EQ_1 = 1.0,
       tsetup_posedge$D$CP$E_EQ_1 = 1.0,
       thold_posedge$D$CP$E_EQ_1 = 1.0,
       tsetup_posedge$E$CP$D_EQ_0 = 1.0,
       thold_posedge$E$CP$D_EQ_0 = 1.0,
       tsetup_posedge$E$CP$D_EQ_1 = 1.0,
       thold_posedge$E$CP$D_EQ_1 = 1.0;

     // path delays
     (posedge CP *> (QN -: E?D:N_S_XM3_G)) = (tpllh$CP$QN, tplhl$CP$QN);
     (posedge CP *> (Q +: E?D:N_S_XM3_G)) = (tpllh$CP$Q, tplhl$CP$Q);
     $setuphold(posedge CP &&& E == 1'b1, negedge D, tsetup_negedge$D$CP$E_EQ_1, thold_negedge$D$CP$E_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& D == 1'b0, negedge E, tsetup_negedge$E$CP$D_EQ_0, thold_negedge$E$CP$D_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& D == 1'b1, negedge E, tsetup_negedge$E$CP$D_EQ_1, thold_negedge$E$CP$D_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& E == 1'b1, posedge D, tsetup_posedge$D$CP$E_EQ_1, thold_posedge$D$CP$E_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& D == 1'b0, posedge E, tsetup_posedge$E$CP$D_EQ_0, thold_posedge$E$CP$D_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& D == 1'b1, posedge E, tsetup_posedge$E$CP$D_EQ_1, thold_posedge$E$CP$D_EQ_1, NOTIFIER);
     $width(posedge CP &&& D_EQ_0_AN_E_EQ_1 == 1'b1, tminpwh$CP$D_EQ_0_AN_E_EQ_1, 0, NOTIFIER);
     $width(negedge CP &&& D_EQ_0_AN_E_EQ_1 == 1'b1, tminpwl$CP$D_EQ_0_AN_E_EQ_1, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF01EHD1 (Q, CP, D, E);
input  CP ;
input  D ;
input  E ;
output Q ;
reg NOTIFIER ;

   udp_mux2 (I0_D, N_S_XM3_G, D, E);
   udp_dff (N_S_XM3_G, I0_D, CP, 1'B0, 1'B0, NOTIFIER);
   not (N_NET0235_XM29_G, N_S_XM3_G);
   not (Q, N_NET0235_XM29_G);
   not (I5_out, D);
   and (D_EQ_0_AN_E_EQ_1, I5_out, E);

   specify
     // delay parameters
     specparam
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tminpwh$CP$D_EQ_0_AN_E_EQ_1 = 1.0,
       tminpwl$CP$D_EQ_0_AN_E_EQ_1 = 1.0,
       tsetup_negedge$D$CP$E_EQ_1 = 1.0,
       thold_negedge$D$CP$E_EQ_1 = 1.0,
       tsetup_negedge$E$CP$D_EQ_0 = 1.0,
       thold_negedge$E$CP$D_EQ_0 = 1.0,
       tsetup_negedge$E$CP$D_EQ_1 = 1.0,
       thold_negedge$E$CP$D_EQ_1 = 1.0,
       tsetup_posedge$D$CP$E_EQ_1 = 1.0,
       thold_posedge$D$CP$E_EQ_1 = 1.0,
       tsetup_posedge$E$CP$D_EQ_0 = 1.0,
       thold_posedge$E$CP$D_EQ_0 = 1.0,
       tsetup_posedge$E$CP$D_EQ_1 = 1.0,
       thold_posedge$E$CP$D_EQ_1 = 1.0;

     // path delays
     (posedge CP *> (Q +: E?D:N_S_XM3_G)) = (tpllh$CP$Q, tplhl$CP$Q);
     $setuphold(posedge CP &&& E == 1'b1, negedge D, tsetup_negedge$D$CP$E_EQ_1, thold_negedge$D$CP$E_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& D == 1'b0, negedge E, tsetup_negedge$E$CP$D_EQ_0, thold_negedge$E$CP$D_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& D == 1'b1, negedge E, tsetup_negedge$E$CP$D_EQ_1, thold_negedge$E$CP$D_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& E == 1'b1, posedge D, tsetup_posedge$D$CP$E_EQ_1, thold_posedge$D$CP$E_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& D == 1'b0, posedge E, tsetup_posedge$E$CP$D_EQ_0, thold_posedge$E$CP$D_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& D == 1'b1, posedge E, tsetup_posedge$E$CP$D_EQ_1, thold_posedge$E$CP$D_EQ_1, NOTIFIER);
     $width(posedge CP &&& D_EQ_0_AN_E_EQ_1 == 1'b1, tminpwh$CP$D_EQ_0_AN_E_EQ_1, 0, NOTIFIER);
     $width(negedge CP &&& D_EQ_0_AN_E_EQ_1 == 1'b1, tminpwl$CP$D_EQ_0_AN_E_EQ_1, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF01EHD2 (Q, CP, D, E);
input  CP ;
input  D ;
input  E ;
output Q ;
reg NOTIFIER ;

   udp_mux2 (I0_D, N_S_XM3_G, D, E);
   udp_dff (N_S_XM3_G, I0_D, CP, 1'B0, 1'B0, NOTIFIER);
   not (N_NET0235_XM29_G, N_S_XM3_G);
   not (Q, N_NET0235_XM29_G);
   not (I5_out, D);
   and (D_EQ_0_AN_E_EQ_1, I5_out, E);

   specify
     // delay parameters
     specparam
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tminpwh$CP$D_EQ_0_AN_E_EQ_1 = 1.0,
       tminpwl$CP$D_EQ_0_AN_E_EQ_1 = 1.0,
       tsetup_negedge$D$CP$E_EQ_1 = 1.0,
       thold_negedge$D$CP$E_EQ_1 = 1.0,
       tsetup_negedge$E$CP$D_EQ_0 = 1.0,
       thold_negedge$E$CP$D_EQ_0 = 1.0,
       tsetup_negedge$E$CP$D_EQ_1 = 1.0,
       thold_negedge$E$CP$D_EQ_1 = 1.0,
       tsetup_posedge$D$CP$E_EQ_1 = 1.0,
       thold_posedge$D$CP$E_EQ_1 = 1.0,
       tsetup_posedge$E$CP$D_EQ_0 = 1.0,
       thold_posedge$E$CP$D_EQ_0 = 1.0,
       tsetup_posedge$E$CP$D_EQ_1 = 1.0,
       thold_posedge$E$CP$D_EQ_1 = 1.0;

     // path delays
     (posedge CP *> (Q +: E?D:N_S_XM3_G)) = (tpllh$CP$Q, tplhl$CP$Q);
     $setuphold(posedge CP &&& E == 1'b1, negedge D, tsetup_negedge$D$CP$E_EQ_1, thold_negedge$D$CP$E_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& D == 1'b0, negedge E, tsetup_negedge$E$CP$D_EQ_0, thold_negedge$E$CP$D_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& D == 1'b1, negedge E, tsetup_negedge$E$CP$D_EQ_1, thold_negedge$E$CP$D_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& E == 1'b1, posedge D, tsetup_posedge$D$CP$E_EQ_1, thold_posedge$D$CP$E_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& D == 1'b0, posedge E, tsetup_posedge$E$CP$D_EQ_0, thold_posedge$E$CP$D_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& D == 1'b1, posedge E, tsetup_posedge$E$CP$D_EQ_1, thold_posedge$E$CP$D_EQ_1, NOTIFIER);
     $width(posedge CP &&& D_EQ_0_AN_E_EQ_1 == 1'b1, tminpwh$CP$D_EQ_0_AN_E_EQ_1, 0, NOTIFIER);
     $width(negedge CP &&& D_EQ_0_AN_E_EQ_1 == 1'b1, tminpwl$CP$D_EQ_0_AN_E_EQ_1, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF01EHD4 (Q, CP, D, E);
input  CP ;
input  D ;
input  E ;
output Q ;
reg NOTIFIER ;

   udp_mux2 (I0_D, N_S_XM3_G, D, E);
   udp_dff (N_S_XM3_G, I0_D, CP, 1'B0, 1'B0, NOTIFIER);
   not (N_NET0235_XM29_G, N_S_XM3_G);
   not (Q, N_NET0235_XM29_G);
   not (I5_out, D);
   and (D_EQ_0_AN_E_EQ_1, I5_out, E);

   specify
     // delay parameters
     specparam
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tminpwh$CP$D_EQ_0_AN_E_EQ_1 = 1.0,
       tminpwl$CP$D_EQ_0_AN_E_EQ_1 = 1.0,
       tsetup_negedge$D$CP$E_EQ_1 = 1.0,
       thold_negedge$D$CP$E_EQ_1 = 1.0,
       tsetup_negedge$E$CP$D_EQ_0 = 1.0,
       thold_negedge$E$CP$D_EQ_0 = 1.0,
       tsetup_negedge$E$CP$D_EQ_1 = 1.0,
       thold_negedge$E$CP$D_EQ_1 = 1.0,
       tsetup_posedge$D$CP$E_EQ_1 = 1.0,
       thold_posedge$D$CP$E_EQ_1 = 1.0,
       tsetup_posedge$E$CP$D_EQ_0 = 1.0,
       thold_posedge$E$CP$D_EQ_0 = 1.0,
       tsetup_posedge$E$CP$D_EQ_1 = 1.0,
       thold_posedge$E$CP$D_EQ_1 = 1.0;

     // path delays
     (posedge CP *> (Q +: E?D:N_S_XM3_G)) = (tpllh$CP$Q, tplhl$CP$Q);
     $setuphold(posedge CP &&& E == 1'b1, negedge D, tsetup_negedge$D$CP$E_EQ_1, thold_negedge$D$CP$E_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& D == 1'b0, negedge E, tsetup_negedge$E$CP$D_EQ_0, thold_negedge$E$CP$D_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& D == 1'b1, negedge E, tsetup_negedge$E$CP$D_EQ_1, thold_negedge$E$CP$D_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& E == 1'b1, posedge D, tsetup_posedge$D$CP$E_EQ_1, thold_posedge$D$CP$E_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& D == 1'b0, posedge E, tsetup_posedge$E$CP$D_EQ_0, thold_posedge$E$CP$D_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& D == 1'b1, posedge E, tsetup_posedge$E$CP$D_EQ_1, thold_posedge$E$CP$D_EQ_1, NOTIFIER);
     $width(posedge CP &&& D_EQ_0_AN_E_EQ_1 == 1'b1, tminpwh$CP$D_EQ_0_AN_E_EQ_1, 0, NOTIFIER);
     $width(negedge CP &&& D_EQ_0_AN_E_EQ_1 == 1'b1, tminpwl$CP$D_EQ_0_AN_E_EQ_1, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF01HD1 (Q, CP, D);
input  CP ;
input  D ;
output Q ;
reg NOTIFIER ;
reg ReSeT;


  
`ifdef  RSTn_lib
	 initial begin
		ReSeT = 0 ;
		#3 ReSeT = 1 ;
		#111 ReSeT = 0 ;
	end

  `else initial  ReSeT = 0;

`endif
 udp_dff (N_S_XM19_G, D, CP, ReSeT , 1'B0, NOTIFIER);

   not (N_NET0130_XM16_D, N_S_XM19_G);
   buf (Q, N_S_XM19_G);

   specify
     // delay parameters
     specparam
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tminpwh$CP$D_EQ_0 = 1.0,
       tminpwl$CP$D_EQ_0 = 1.0,
       tsetup_negedge$D$CP = 1.0,
       thold_negedge$D$CP = 1.0,
       tsetup_posedge$D$CP = 1.0,
       thold_posedge$D$CP = 1.0;

     // path delays
     (posedge CP *> (Q +: D)) = (tpllh$CP$Q, tplhl$CP$Q);
     $setuphold(posedge CP, negedge D, tsetup_negedge$D$CP, thold_negedge$D$CP, NOTIFIER);
     $setuphold(posedge CP, posedge D, tsetup_posedge$D$CP, thold_posedge$D$CP, NOTIFIER);
     $width(posedge CP &&& D == 1'b0, tminpwh$CP$D_EQ_0, 0, NOTIFIER);
     $width(negedge CP &&& D == 1'b0, tminpwl$CP$D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF01HD2 (Q, CP, D);
input  CP ;
input  D ;
output Q ;
reg NOTIFIER ;

reg ReSeT;

 
 `ifdef  RSTn_lib
	 initial begin
		ReSeT = 0 ;
		#3 ReSeT = 1 ;
		#111 ReSeT = 0 ;
	end

  `else initial  ReSeT = 0;

`endif
   udp_dff (N_S_XM19_G, D, CP, ReSeT, 1'B0, NOTIFIER);
 not (N_NET0130_XM16_D, N_S_XM19_G);
   buf (Q, N_S_XM19_G);

   specify
     // delay parameters
     specparam
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tminpwh$CP$D_EQ_0 = 1.0,
       tminpwl$CP$D_EQ_0 = 1.0,
       tsetup_negedge$D$CP = 1.0,
       thold_negedge$D$CP = 1.0,
       tsetup_posedge$D$CP = 1.0,
       thold_posedge$D$CP = 1.0;

     // path delays
     (posedge CP *> (Q +: D)) = (tpllh$CP$Q, tplhl$CP$Q);
     $setuphold(posedge CP, negedge D, tsetup_negedge$D$CP, thold_negedge$D$CP, NOTIFIER);
     $setuphold(posedge CP, posedge D, tsetup_posedge$D$CP, thold_posedge$D$CP, NOTIFIER);
     $width(posedge CP &&& D == 1'b0, tminpwh$CP$D_EQ_0, 0, NOTIFIER);
     $width(negedge CP &&& D == 1'b0, tminpwl$CP$D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF01HD4 (Q, CP, D);
input  CP ;
input  D ;
output Q ;
reg NOTIFIER ;
reg ReSeT;


`ifdef  RSTn_lib
	 initial begin
		ReSeT = 0 ;
		#3 ReSeT = 1 ;
		#111 ReSeT = 0 ;
	end
  `else initial  ReSeT = 0;
`endif
   udp_dff (N_S_XM19_G, D, CP, ReSeT , 1'B0, NOTIFIER);
   not (N_NET0130_XM16_D, N_S_XM19_G);
   buf (Q, N_S_XM19_G);

   specify
     // delay parameters
     specparam
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tminpwh$CP$D_EQ_0 = 1.0,
       tminpwl$CP$D_EQ_0 = 1.0,
       tsetup_negedge$D$CP = 1.0,
       thold_negedge$D$CP = 1.0,
       tsetup_posedge$D$CP = 1.0,
       thold_posedge$D$CP = 1.0;

     // path delays
     (posedge CP *> (Q +: D)) = (tpllh$CP$Q, tplhl$CP$Q);
     $setuphold(posedge CP, negedge D, tsetup_negedge$D$CP, thold_negedge$D$CP, NOTIFIER);
     $setuphold(posedge CP, posedge D, tsetup_posedge$D$CP, thold_posedge$D$CP, NOTIFIER);
     $width(posedge CP &&& D == 1'b0, tminpwh$CP$D_EQ_0, 0, NOTIFIER);
     $width(negedge CP &&& D == 1'b0, tminpwl$CP$D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF02D1 (Q, QN, CDN, CP, D);
input  CDN ;
input  CP ;
input  D ;
output Q ;
output QN ;
reg NOTIFIER ;

   not (I0_CLEAR, CDN);
   udp_dff (N_S_XM23_G, D, CP, I0_CLEAR, 1'B0, NOTIFIER);
   not (N_NET0130_XM20_D, N_S_XM23_G);
   buf (Q, N_S_XM23_G);
   not (QN, N_S_XM23_G);
   not (I7_out, D);
   and (CDN_EQ_1_AN_D_EQ_0, CDN, I7_out);

   specify
     // delay parameters
     specparam
       tphhl$CDN$Q = 1.0,
       tphlh$CDN$QN = 1.0,
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tpllh$CP$QN = 1.0,
       tplhl$CP$QN = 1.0,
       tminpwl$CDN$D_EQ_0 = 1.0,
       tminpwh$CP$CDN_EQ_1_AN_D_EQ_0 = 1.0,
       tminpwl$CP$CDN_EQ_1_AN_D_EQ_0 = 1.0,
       tsetup_negedge$D$CP$CDN_EQ_1 = 1.0,
       thold_negedge$D$CP$CDN_EQ_1 = 1.0,
       tsetup_posedge$D$CP$CDN_EQ_1 = 1.0,
       thold_posedge$D$CP$CDN_EQ_1 = 1.0,
       trec$CDN$CP$D_EQ_1 = 1.0,
       trem$CDN$CP$D_EQ_1 = 1.0;

     // path delays
     (posedge CP *> (QN -: D)) = (tpllh$CP$QN, tplhl$CP$QN);
     (posedge CP *> (Q +: D)) = (tpllh$CP$Q, tplhl$CP$Q);
     (negedge CDN *> (QN +: 1'b1)) = (tphlh$CDN$QN, 0);
     (negedge CDN *> (Q -: 1'b1)) = (0, tphhl$CDN$Q);
     $setuphold(posedge CP &&& CDN == 1'b1, negedge D, tsetup_negedge$D$CP$CDN_EQ_1, thold_negedge$D$CP$CDN_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& CDN == 1'b1, posedge D, tsetup_posedge$D$CP$CDN_EQ_1, thold_posedge$D$CP$CDN_EQ_1, NOTIFIER);
     $recrem(posedge CDN, posedge CP &&& D == 1'b1, trec$CDN$CP$D_EQ_1, trem$CDN$CP$D_EQ_1, NOTIFIER);
     $width(negedge CDN &&& D == 1'b0, tminpwl$CDN$D_EQ_0, 0, NOTIFIER);
     $width(posedge CP &&& CDN_EQ_1_AN_D_EQ_0 == 1'b1, tminpwh$CP$CDN_EQ_1_AN_D_EQ_0, 0, NOTIFIER);
     $width(negedge CP &&& CDN_EQ_1_AN_D_EQ_0 == 1'b1, tminpwl$CP$CDN_EQ_1_AN_D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF02D2 (Q, QN, CDN, CP, D);
input  CDN ;
input  CP ;
input  D ;
output Q ;
output QN ;
reg NOTIFIER ;

   not (I0_CLEAR, CDN);
   udp_dff (N_S_XM23_G, D, CP, I0_CLEAR, 1'B0, NOTIFIER);
   not (N_NET0130_XM20_D, N_S_XM23_G);
   buf (Q, N_S_XM23_G);
   not (QN, N_S_XM23_G);
   not (I7_out, D);
   and (CDN_EQ_1_AN_D_EQ_0, CDN, I7_out);

   specify
     // delay parameters
     specparam
       tphhl$CDN$Q = 1.0,
       tphlh$CDN$QN = 1.0,
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tpllh$CP$QN = 1.0,
       tplhl$CP$QN = 1.0,
       tminpwl$CDN$D_EQ_0 = 1.0,
       tminpwh$CP$CDN_EQ_1_AN_D_EQ_0 = 1.0,
       tminpwl$CP$CDN_EQ_1_AN_D_EQ_0 = 1.0,
       tsetup_negedge$D$CP$CDN_EQ_1 = 1.0,
       thold_negedge$D$CP$CDN_EQ_1 = 1.0,
       tsetup_posedge$D$CP$CDN_EQ_1 = 1.0,
       thold_posedge$D$CP$CDN_EQ_1 = 1.0,
       trec$CDN$CP$D_EQ_1 = 1.0,
       trem$CDN$CP$D_EQ_1 = 1.0;

     // path delays
     (posedge CP *> (QN -: D)) = (tpllh$CP$QN, tplhl$CP$QN);
     (posedge CP *> (Q +: D)) = (tpllh$CP$Q, tplhl$CP$Q);
     (negedge CDN *> (QN +: 1'b1)) = (tphlh$CDN$QN, 0);
     (negedge CDN *> (Q -: 1'b1)) = (0, tphhl$CDN$Q);
     $setuphold(posedge CP &&& CDN == 1'b1, negedge D, tsetup_negedge$D$CP$CDN_EQ_1, thold_negedge$D$CP$CDN_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& CDN == 1'b1, posedge D, tsetup_posedge$D$CP$CDN_EQ_1, thold_posedge$D$CP$CDN_EQ_1, NOTIFIER);
     $recrem(posedge CDN, posedge CP &&& D == 1'b1, trec$CDN$CP$D_EQ_1, trem$CDN$CP$D_EQ_1, NOTIFIER);
     $width(negedge CDN &&& D == 1'b0, tminpwl$CDN$D_EQ_0, 0, NOTIFIER);
     $width(posedge CP &&& CDN_EQ_1_AN_D_EQ_0 == 1'b1, tminpwh$CP$CDN_EQ_1_AN_D_EQ_0, 0, NOTIFIER);
     $width(negedge CP &&& CDN_EQ_1_AN_D_EQ_0 == 1'b1, tminpwl$CP$CDN_EQ_1_AN_D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF02D4 (Q, QN, CDN, CP, D);
input  CDN ;
input  CP ;
input  D ;
output Q ;
output QN ;
reg NOTIFIER ;

   not (I0_CLEAR, CDN);
   udp_dff (N_S_XM23_G, D, CP, I0_CLEAR, 1'B0, NOTIFIER);
   not (N_NET0130_XM20_D, N_S_XM23_G);
   buf (Q, N_S_XM23_G);
   not (QN, N_S_XM23_G);
   not (I7_out, D);
   and (CDN_EQ_1_AN_D_EQ_0, CDN, I7_out);

   specify
     // delay parameters
     specparam
       tphhl$CDN$Q = 1.0,
       tphlh$CDN$QN = 1.0,
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tpllh$CP$QN = 1.0,
       tplhl$CP$QN = 1.0,
       tminpwl$CDN$D_EQ_0 = 1.0,
       tminpwh$CP$CDN_EQ_1_AN_D_EQ_0 = 1.0,
       tminpwl$CP$CDN_EQ_1_AN_D_EQ_0 = 1.0,
       tsetup_negedge$D$CP$CDN_EQ_1 = 1.0,
       thold_negedge$D$CP$CDN_EQ_1 = 1.0,
       tsetup_posedge$D$CP$CDN_EQ_1 = 1.0,
       thold_posedge$D$CP$CDN_EQ_1 = 1.0,
       trec$CDN$CP$D_EQ_1 = 1.0,
       trem$CDN$CP$D_EQ_1 = 1.0;

     // path delays
     (posedge CP *> (QN -: D)) = (tpllh$CP$QN, tplhl$CP$QN);
     (posedge CP *> (Q +: D)) = (tpllh$CP$Q, tplhl$CP$Q);
     (negedge CDN *> (QN +: 1'b1)) = (tphlh$CDN$QN, 0);
     (negedge CDN *> (Q -: 1'b1)) = (0, tphhl$CDN$Q);
     $setuphold(posedge CP &&& CDN == 1'b1, negedge D, tsetup_negedge$D$CP$CDN_EQ_1, thold_negedge$D$CP$CDN_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& CDN == 1'b1, posedge D, tsetup_posedge$D$CP$CDN_EQ_1, thold_posedge$D$CP$CDN_EQ_1, NOTIFIER);
     $recrem(posedge CDN, posedge CP &&& D == 1'b1, trec$CDN$CP$D_EQ_1, trem$CDN$CP$D_EQ_1, NOTIFIER);
     $width(negedge CDN &&& D == 1'b0, tminpwl$CDN$D_EQ_0, 0, NOTIFIER);
     $width(posedge CP &&& CDN_EQ_1_AN_D_EQ_0 == 1'b1, tminpwh$CP$CDN_EQ_1_AN_D_EQ_0, 0, NOTIFIER);
     $width(negedge CP &&& CDN_EQ_1_AN_D_EQ_0 == 1'b1, tminpwl$CP$CDN_EQ_1_AN_D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF02ED1 (Q, QN, CDN, CP, D, E);
input  CDN ;
input  CP ;
input  D ;
input  E ;
output Q ;
output QN ;
reg NOTIFIER ;

   udp_mux2 (I0_D, N_S_XM3_G, D, E);
   not (I0_CLEAR, CDN);
   udp_dff (N_S_XM3_G, I0_D, CP, I0_CLEAR, 1'B0, NOTIFIER);
   not (N_NET0235_XM31_G, N_S_XM3_G);
   not (Q, N_NET0235_XM31_G);
   not (QN, N_S_XM3_G);
   and (CDN_EQ_1_AN_E_EQ_1, CDN, E);
   and (D_EQ_1_AN_E_EQ_1, D, E);
   not (I9_out, D);
   not (I10_out, E);
   and (D_EQ_0_AN_E_EQ_0, I9_out, I10_out);
   not (I12_out, D);
   and (CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1, CDN, I12_out, E);

   specify
     // delay parameters
     specparam
       tphhl$CDN$Q = 1.0,
       tphlh$CDN$QN = 1.0,
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tpllh$CP$QN = 1.0,
       tplhl$CP$QN = 1.0,
       tminpwl$CDN$D_EQ_0_AN_E_EQ_0 = 1.0,
       tminpwh$CP$CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1 = 1.0,
       tminpwl$CP$CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1 = 1.0,
       tsetup_negedge$D$CP$CDN_EQ_1_AN_E_EQ_1 = 1.0,
       thold_negedge$D$CP$CDN_EQ_1_AN_E_EQ_1 = 1.0,
       tsetup_negedge$E$CP$CDN_EQ_1 = 1.0,
       thold_negedge$E$CP$CDN_EQ_1 = 1.0,
       tsetup_posedge$D$CP$CDN_EQ_1_AN_E_EQ_1 = 1.0,
       thold_posedge$D$CP$CDN_EQ_1_AN_E_EQ_1 = 1.0,
       tsetup_posedge$E$CP$CDN_EQ_1 = 1.0,
       thold_posedge$E$CP$CDN_EQ_1 = 1.0,
       trec$CDN$CP$D_EQ_1_AN_E_EQ_1 = 1.0,
       trem$CDN$CP$D_EQ_1_AN_E_EQ_1 = 1.0;

     // path delays
     (posedge CP *> (QN -: E?D:N_S_XM3_G)) = (tpllh$CP$QN, tplhl$CP$QN);
     (posedge CP *> (Q +: E?D:N_S_XM3_G)) = (tpllh$CP$Q, tplhl$CP$Q);
     (negedge CDN *> (QN +: 1'b1)) = (tphlh$CDN$QN, 0);
     (negedge CDN *> (Q -: 1'b1)) = (0, tphhl$CDN$Q);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_E_EQ_1 == 1'b1, negedge D, tsetup_negedge$D$CP$CDN_EQ_1_AN_E_EQ_1, thold_negedge$D$CP$CDN_EQ_1_AN_E_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& CDN == 1'b1, negedge E, tsetup_negedge$E$CP$CDN_EQ_1, thold_negedge$E$CP$CDN_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_E_EQ_1 == 1'b1, posedge D, tsetup_posedge$D$CP$CDN_EQ_1_AN_E_EQ_1, thold_posedge$D$CP$CDN_EQ_1_AN_E_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& CDN == 1'b1, posedge E, tsetup_posedge$E$CP$CDN_EQ_1, thold_posedge$E$CP$CDN_EQ_1, NOTIFIER);
     $recrem(posedge CDN, posedge CP &&& D_EQ_1_AN_E_EQ_1 == 1'b1, trec$CDN$CP$D_EQ_1_AN_E_EQ_1, trem$CDN$CP$D_EQ_1_AN_E_EQ_1, NOTIFIER);
     $width(negedge CDN &&& D_EQ_0_AN_E_EQ_0 == 1'b1, tminpwl$CDN$D_EQ_0_AN_E_EQ_0, 0, NOTIFIER);
     $width(posedge CP &&& CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1 == 1'b1, tminpwh$CP$CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1, 0, NOTIFIER);
     $width(negedge CP &&& CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1 == 1'b1, tminpwl$CP$CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF02ED2 (Q, QN, CDN, CP, D, E);
input  CDN ;
input  CP ;
input  D ;
input  E ;
output Q ;
output QN ;
reg NOTIFIER ;

   udp_mux2 (I0_D, N_S_XM3_G, D, E);
   not (I0_CLEAR, CDN);
   udp_dff (N_S_XM3_G, I0_D, CP, I0_CLEAR, 1'B0, NOTIFIER);
   not (N_NET0235_XM31_G, N_S_XM3_G);
   not (Q, N_NET0235_XM31_G);
   not (QN, N_S_XM3_G);
   and (CDN_EQ_1_AN_E_EQ_1, CDN, E);
   and (D_EQ_1_AN_E_EQ_1, D, E);
   not (I9_out, D);
   not (I10_out, E);
   and (D_EQ_0_AN_E_EQ_0, I9_out, I10_out);
   not (I12_out, D);
   and (CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1, CDN, I12_out, E);

   specify
     // delay parameters
     specparam
       tphhl$CDN$Q = 1.0,
       tphlh$CDN$QN = 1.0,
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tpllh$CP$QN = 1.0,
       tplhl$CP$QN = 1.0,
       tminpwl$CDN$D_EQ_0_AN_E_EQ_0 = 1.0,
       tminpwh$CP$CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1 = 1.0,
       tminpwl$CP$CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1 = 1.0,
       tsetup_negedge$D$CP$CDN_EQ_1_AN_E_EQ_1 = 1.0,
       thold_negedge$D$CP$CDN_EQ_1_AN_E_EQ_1 = 1.0,
       tsetup_negedge$E$CP$CDN_EQ_1 = 1.0,
       thold_negedge$E$CP$CDN_EQ_1 = 1.0,
       tsetup_posedge$D$CP$CDN_EQ_1_AN_E_EQ_1 = 1.0,
       thold_posedge$D$CP$CDN_EQ_1_AN_E_EQ_1 = 1.0,
       tsetup_posedge$E$CP$CDN_EQ_1 = 1.0,
       thold_posedge$E$CP$CDN_EQ_1 = 1.0,
       trec$CDN$CP$D_EQ_1_AN_E_EQ_1 = 1.0,
       trem$CDN$CP$D_EQ_1_AN_E_EQ_1 = 1.0;

     // path delays
     (posedge CP *> (QN -: E?D:N_S_XM3_G)) = (tpllh$CP$QN, tplhl$CP$QN);
     (posedge CP *> (Q +: E?D:N_S_XM3_G)) = (tpllh$CP$Q, tplhl$CP$Q);
     (negedge CDN *> (QN +: 1'b1)) = (tphlh$CDN$QN, 0);
     (negedge CDN *> (Q -: 1'b1)) = (0, tphhl$CDN$Q);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_E_EQ_1 == 1'b1, negedge D, tsetup_negedge$D$CP$CDN_EQ_1_AN_E_EQ_1, thold_negedge$D$CP$CDN_EQ_1_AN_E_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& CDN == 1'b1, negedge E, tsetup_negedge$E$CP$CDN_EQ_1, thold_negedge$E$CP$CDN_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_E_EQ_1 == 1'b1, posedge D, tsetup_posedge$D$CP$CDN_EQ_1_AN_E_EQ_1, thold_posedge$D$CP$CDN_EQ_1_AN_E_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& CDN == 1'b1, posedge E, tsetup_posedge$E$CP$CDN_EQ_1, thold_posedge$E$CP$CDN_EQ_1, NOTIFIER);
     $recrem(posedge CDN, posedge CP &&& D_EQ_1_AN_E_EQ_1 == 1'b1, trec$CDN$CP$D_EQ_1_AN_E_EQ_1, trem$CDN$CP$D_EQ_1_AN_E_EQ_1, NOTIFIER);
     $width(negedge CDN &&& D_EQ_0_AN_E_EQ_0 == 1'b1, tminpwl$CDN$D_EQ_0_AN_E_EQ_0, 0, NOTIFIER);
     $width(posedge CP &&& CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1 == 1'b1, tminpwh$CP$CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1, 0, NOTIFIER);
     $width(negedge CP &&& CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1 == 1'b1, tminpwl$CP$CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF02ED4 (Q, QN, CDN, CP, D, E);
input  CDN ;
input  CP ;
input  D ;
input  E ;
output Q ;
output QN ;
reg NOTIFIER ;

   udp_mux2 (I0_D, N_S_XM3_G, D, E);
   not (I0_CLEAR, CDN);
   udp_dff (N_S_XM3_G, I0_D, CP, I0_CLEAR, 1'B0, NOTIFIER);
   not (N_NET0235_XM31_G, N_S_XM3_G);
   not (Q, N_NET0235_XM31_G);
   not (QN, N_S_XM3_G);
   and (CDN_EQ_1_AN_E_EQ_1, CDN, E);
   and (D_EQ_1_AN_E_EQ_1, D, E);
   not (I9_out, D);
   not (I10_out, E);
   and (D_EQ_0_AN_E_EQ_0, I9_out, I10_out);
   not (I12_out, D);
   and (CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1, CDN, I12_out, E);

   specify
     // delay parameters
     specparam
       tphhl$CDN$Q = 1.0,
       tphlh$CDN$QN = 1.0,
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tpllh$CP$QN = 1.0,
       tplhl$CP$QN = 1.0,
       tminpwl$CDN$D_EQ_0_AN_E_EQ_0 = 1.0,
       tminpwh$CP$CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1 = 1.0,
       tminpwl$CP$CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1 = 1.0,
       tsetup_negedge$D$CP$CDN_EQ_1_AN_E_EQ_1 = 1.0,
       thold_negedge$D$CP$CDN_EQ_1_AN_E_EQ_1 = 1.0,
       tsetup_negedge$E$CP$CDN_EQ_1 = 1.0,
       thold_negedge$E$CP$CDN_EQ_1 = 1.0,
       tsetup_posedge$D$CP$CDN_EQ_1_AN_E_EQ_1 = 1.0,
       thold_posedge$D$CP$CDN_EQ_1_AN_E_EQ_1 = 1.0,
       tsetup_posedge$E$CP$CDN_EQ_1 = 1.0,
       thold_posedge$E$CP$CDN_EQ_1 = 1.0,
       trec$CDN$CP$D_EQ_1_AN_E_EQ_1 = 1.0,
       trem$CDN$CP$D_EQ_1_AN_E_EQ_1 = 1.0;

     // path delays
     (posedge CP *> (QN -: E?D:N_S_XM3_G)) = (tpllh$CP$QN, tplhl$CP$QN);
     (posedge CP *> (Q +: E?D:N_S_XM3_G)) = (tpllh$CP$Q, tplhl$CP$Q);
     (negedge CDN *> (QN +: 1'b1)) = (tphlh$CDN$QN, 0);
     (negedge CDN *> (Q -: 1'b1)) = (0, tphhl$CDN$Q);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_E_EQ_1 == 1'b1, negedge D, tsetup_negedge$D$CP$CDN_EQ_1_AN_E_EQ_1, thold_negedge$D$CP$CDN_EQ_1_AN_E_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& CDN == 1'b1, negedge E, tsetup_negedge$E$CP$CDN_EQ_1, thold_negedge$E$CP$CDN_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_E_EQ_1 == 1'b1, posedge D, tsetup_posedge$D$CP$CDN_EQ_1_AN_E_EQ_1, thold_posedge$D$CP$CDN_EQ_1_AN_E_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& CDN == 1'b1, posedge E, tsetup_posedge$E$CP$CDN_EQ_1, thold_posedge$E$CP$CDN_EQ_1, NOTIFIER);
     $recrem(posedge CDN, posedge CP &&& D_EQ_1_AN_E_EQ_1 == 1'b1, trec$CDN$CP$D_EQ_1_AN_E_EQ_1, trem$CDN$CP$D_EQ_1_AN_E_EQ_1, NOTIFIER);
     $width(negedge CDN &&& D_EQ_0_AN_E_EQ_0 == 1'b1, tminpwl$CDN$D_EQ_0_AN_E_EQ_0, 0, NOTIFIER);
     $width(posedge CP &&& CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1 == 1'b1, tminpwh$CP$CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1, 0, NOTIFIER);
     $width(negedge CP &&& CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1 == 1'b1, tminpwl$CP$CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF02HD1 (Q, CDN, CP, D);
input  CDN ;
input  CP ;
input  D ;
output Q ;
reg NOTIFIER ;

   not (I0_CLEAR, CDN);
   udp_dff (N_S_XM23_G, D, CP, I0_CLEAR, 1'B0, NOTIFIER);
   not (N_NET0130_XM20_D, N_S_XM23_G);
   not (Q, N_NET0130_XM20_D);
   not (I5_out, D);
   and (CDN_EQ_1_AN_D_EQ_0, CDN, I5_out);

   specify
     // delay parameters
     specparam
       tphhl$CDN$Q = 1.0,
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tminpwl$CDN$D_EQ_0 = 1.0,
       tminpwh$CP$CDN_EQ_1_AN_D_EQ_0 = 1.0,
       tminpwl$CP$CDN_EQ_1_AN_D_EQ_0 = 1.0,
       tsetup_negedge$D$CP$CDN_EQ_1 = 1.0,
       thold_negedge$D$CP$CDN_EQ_1 = 1.0,
       tsetup_posedge$D$CP$CDN_EQ_1 = 1.0,
       thold_posedge$D$CP$CDN_EQ_1 = 1.0,
       trec$CDN$CP$D_EQ_1 = 1.0,
       trem$CDN$CP$D_EQ_1 = 1.0;

     // path delays
     (posedge CP *> (Q +: D)) = (tpllh$CP$Q, tplhl$CP$Q);
     (negedge CDN *> (Q -: 1'b1)) = (0, tphhl$CDN$Q);
     $setuphold(posedge CP &&& CDN == 1'b1, negedge D, tsetup_negedge$D$CP$CDN_EQ_1, thold_negedge$D$CP$CDN_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& CDN == 1'b1, posedge D, tsetup_posedge$D$CP$CDN_EQ_1, thold_posedge$D$CP$CDN_EQ_1, NOTIFIER);
     $recrem(posedge CDN, posedge CP &&& D == 1'b1, trec$CDN$CP$D_EQ_1, trem$CDN$CP$D_EQ_1, NOTIFIER);
     $width(negedge CDN &&& D == 1'b0, tminpwl$CDN$D_EQ_0, 0, NOTIFIER);
     $width(posedge CP &&& CDN_EQ_1_AN_D_EQ_0 == 1'b1, tminpwh$CP$CDN_EQ_1_AN_D_EQ_0, 0, NOTIFIER);
     $width(negedge CP &&& CDN_EQ_1_AN_D_EQ_0 == 1'b1, tminpwl$CP$CDN_EQ_1_AN_D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF02HD2 (Q, CDN, CP, D);
input  CDN ;
input  CP ;
input  D ;
output Q ;
reg NOTIFIER ;

   not (I0_CLEAR, CDN);
   udp_dff (N_S_XM23_G, D, CP, I0_CLEAR, 1'B0, NOTIFIER);
   not (N_NET0130_XM20_D, N_S_XM23_G);
   not (Q, N_NET0130_XM20_D);
   not (I5_out, D);
   and (CDN_EQ_1_AN_D_EQ_0, CDN, I5_out);

   specify
     // delay parameters
     specparam
       tphhl$CDN$Q = 1.0,
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tminpwl$CDN$D_EQ_0 = 1.0,
       tminpwh$CP$CDN_EQ_1_AN_D_EQ_0 = 1.0,
       tminpwl$CP$CDN_EQ_1_AN_D_EQ_0 = 1.0,
       tsetup_negedge$D$CP$CDN_EQ_1 = 1.0,
       thold_negedge$D$CP$CDN_EQ_1 = 1.0,
       tsetup_posedge$D$CP$CDN_EQ_1 = 1.0,
       thold_posedge$D$CP$CDN_EQ_1 = 1.0,
       trec$CDN$CP$D_EQ_1 = 1.0,
       trem$CDN$CP$D_EQ_1 = 1.0;

     // path delays
     (posedge CP *> (Q +: D)) = (tpllh$CP$Q, tplhl$CP$Q);
     (negedge CDN *> (Q -: 1'b1)) = (0, tphhl$CDN$Q);
     $setuphold(posedge CP &&& CDN == 1'b1, negedge D, tsetup_negedge$D$CP$CDN_EQ_1, thold_negedge$D$CP$CDN_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& CDN == 1'b1, posedge D, tsetup_posedge$D$CP$CDN_EQ_1, thold_posedge$D$CP$CDN_EQ_1, NOTIFIER);
     $recrem(posedge CDN, posedge CP &&& D == 1'b1, trec$CDN$CP$D_EQ_1, trem$CDN$CP$D_EQ_1, NOTIFIER);
     $width(negedge CDN &&& D == 1'b0, tminpwl$CDN$D_EQ_0, 0, NOTIFIER);
     $width(posedge CP &&& CDN_EQ_1_AN_D_EQ_0 == 1'b1, tminpwh$CP$CDN_EQ_1_AN_D_EQ_0, 0, NOTIFIER);
     $width(negedge CP &&& CDN_EQ_1_AN_D_EQ_0 == 1'b1, tminpwl$CP$CDN_EQ_1_AN_D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF02HD4 (Q, CDN, CP, D);
input  CDN ;
input  CP ;
input  D ;
output Q ;
reg NOTIFIER ;

   not (I0_CLEAR, CDN);
   udp_dff (N_S_XM23_G, D, CP, I0_CLEAR, 1'B0, NOTIFIER);
   not (N_NET0130_XM20_D, N_S_XM23_G);
   not (Q, N_NET0130_XM20_D);
   not (I5_out, D);
   and (CDN_EQ_1_AN_D_EQ_0, CDN, I5_out);

   specify
     // delay parameters
     specparam
       tphhl$CDN$Q = 1.0,
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tminpwl$CDN$D_EQ_0 = 1.0,
       tminpwh$CP$CDN_EQ_1_AN_D_EQ_0 = 1.0,
       tminpwl$CP$CDN_EQ_1_AN_D_EQ_0 = 1.0,
       tsetup_negedge$D$CP$CDN_EQ_1 = 1.0,
       thold_negedge$D$CP$CDN_EQ_1 = 1.0,
       tsetup_posedge$D$CP$CDN_EQ_1 = 1.0,
       thold_posedge$D$CP$CDN_EQ_1 = 1.0,
       trec$CDN$CP$D_EQ_1 = 1.0,
       trem$CDN$CP$D_EQ_1 = 1.0;

     // path delays
     (posedge CP *> (Q +: D)) = (tpllh$CP$Q, tplhl$CP$Q);
     (negedge CDN *> (Q -: 1'b1)) = (0, tphhl$CDN$Q);
     $setuphold(posedge CP &&& CDN == 1'b1, negedge D, tsetup_negedge$D$CP$CDN_EQ_1, thold_negedge$D$CP$CDN_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& CDN == 1'b1, posedge D, tsetup_posedge$D$CP$CDN_EQ_1, thold_posedge$D$CP$CDN_EQ_1, NOTIFIER);
     $recrem(posedge CDN, posedge CP &&& D == 1'b1, trec$CDN$CP$D_EQ_1, trem$CDN$CP$D_EQ_1, NOTIFIER);
     $width(negedge CDN &&& D == 1'b0, tminpwl$CDN$D_EQ_0, 0, NOTIFIER);
     $width(posedge CP &&& CDN_EQ_1_AN_D_EQ_0 == 1'b1, tminpwh$CP$CDN_EQ_1_AN_D_EQ_0, 0, NOTIFIER);
     $width(negedge CP &&& CDN_EQ_1_AN_D_EQ_0 == 1'b1, tminpwl$CP$CDN_EQ_1_AN_D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF03D1 (Q, QN, CP, D, SDN);
input  CP ;
input  D ;
input  SDN ;
output Q ;
output QN ;
reg NOTIFIER ;
reg ReSeT;
`ifdef  RSTn_lib
    
	 initial begin
		ReSeT = 0 ;
		#3 ReSeT = 1 ;
		#111 ReSeT = 0 ;
	end
  `else initial  ReSeT = 0;
`endif

   not (I0_SET, SDN);
   udp_dff (N_S_XM21_G, D, CP, ReSeT , I0_SET, NOTIFIER);


   not (N_NET0130_XM18_D, N_S_XM21_G);
   buf (Q, N_S_XM21_G);
   not (QN, N_S_XM21_G);
   not (I7_out, D);
   and (D_EQ_0_AN_SDN_EQ_1, I7_out, SDN);

   specify
     // delay parameters
     specparam
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tpllh$CP$QN = 1.0,
       tplhl$CP$QN = 1.0,
       tphlh$SDN$Q = 1.0,
       tphhl$SDN$QN = 1.0,
       tminpwh$CP$D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwl$CP$D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwl$SDN$D_EQ_0 = 1.0,
       tsetup_negedge$D$CP$SDN_EQ_1 = 1.0,
       thold_negedge$D$CP$SDN_EQ_1 = 1.0,
       tsetup_posedge$D$CP$SDN_EQ_1 = 1.0,
       thold_posedge$D$CP$SDN_EQ_1 = 1.0,
       trec$SDN$CP$D_EQ_0 = 1.0,
       trem$SDN$CP$D_EQ_0 = 1.0;

     // path delays
     (posedge CP *> (QN -: D)) = (tpllh$CP$QN, tplhl$CP$QN);
     (posedge CP *> (Q +: D)) = (tpllh$CP$Q, tplhl$CP$Q);
     (negedge SDN *> (QN -: 1'b1)) = (0, tphhl$SDN$QN);
     (negedge SDN *> (Q +: 1'b1)) = (tphlh$SDN$Q, 0);
     $setuphold(posedge CP &&& SDN == 1'b1, negedge D, tsetup_negedge$D$CP$SDN_EQ_1, thold_negedge$D$CP$SDN_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& SDN == 1'b1, posedge D, tsetup_posedge$D$CP$SDN_EQ_1, thold_posedge$D$CP$SDN_EQ_1, NOTIFIER);
     $recrem(posedge SDN, posedge CP &&& D == 1'b0, trec$SDN$CP$D_EQ_0, trem$SDN$CP$D_EQ_0, NOTIFIER);
     $width(posedge CP &&& D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwh$CP$D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(negedge CP &&& D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwl$CP$D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(negedge SDN &&& D == 1'b0, tminpwl$SDN$D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF03D2 (Q, QN, CP, D, SDN);
input  CP ;
input  D ;
input  SDN ;
output Q ;
output QN ;
reg NOTIFIER ;

   not (I0_SET, SDN);
   udp_dff (N_S_XM21_G, D, CP, 1'B0, I0_SET, NOTIFIER);
   not (N_NET0130_XM18_D, N_S_XM21_G);
   buf (Q, N_S_XM21_G);
   not (QN, N_S_XM21_G);
   not (I7_out, D);
   and (D_EQ_0_AN_SDN_EQ_1, I7_out, SDN);

   specify
     // delay parameters
     specparam
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tpllh$CP$QN = 1.0,
       tplhl$CP$QN = 1.0,
       tphlh$SDN$Q = 1.0,
       tphhl$SDN$QN = 1.0,
       tminpwh$CP$D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwl$CP$D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwl$SDN$D_EQ_0 = 1.0,
       tsetup_negedge$D$CP$SDN_EQ_1 = 1.0,
       thold_negedge$D$CP$SDN_EQ_1 = 1.0,
       tsetup_posedge$D$CP$SDN_EQ_1 = 1.0,
       thold_posedge$D$CP$SDN_EQ_1 = 1.0,
       trec$SDN$CP$D_EQ_0 = 1.0,
       trem$SDN$CP$D_EQ_0 = 1.0;

     // path delays
     (posedge CP *> (QN -: D)) = (tpllh$CP$QN, tplhl$CP$QN);
     (posedge CP *> (Q +: D)) = (tpllh$CP$Q, tplhl$CP$Q);
     (negedge SDN *> (QN -: 1'b1)) = (0, tphhl$SDN$QN);
     (negedge SDN *> (Q +: 1'b1)) = (tphlh$SDN$Q, 0);
     $setuphold(posedge CP &&& SDN == 1'b1, negedge D, tsetup_negedge$D$CP$SDN_EQ_1, thold_negedge$D$CP$SDN_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& SDN == 1'b1, posedge D, tsetup_posedge$D$CP$SDN_EQ_1, thold_posedge$D$CP$SDN_EQ_1, NOTIFIER);
     $recrem(posedge SDN, posedge CP &&& D == 1'b0, trec$SDN$CP$D_EQ_0, trem$SDN$CP$D_EQ_0, NOTIFIER);
     $width(posedge CP &&& D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwh$CP$D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(negedge CP &&& D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwl$CP$D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(negedge SDN &&& D == 1'b0, tminpwl$SDN$D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF03D4 (Q, QN, CP, D, SDN);
input  CP ;
input  D ;
input  SDN ;
output Q ;
output QN ;
reg NOTIFIER ;

   not (I0_SET, SDN);
   udp_dff (N_S_XM21_G, D, CP, 1'B0, I0_SET, NOTIFIER);
   not (N_NET0130_XM18_D, N_S_XM21_G);
   buf (Q, N_S_XM21_G);
   not (QN, N_S_XM21_G);
   not (I7_out, D);
   and (D_EQ_0_AN_SDN_EQ_1, I7_out, SDN);

   specify
     // delay parameters
     specparam
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tpllh$CP$QN = 1.0,
       tplhl$CP$QN = 1.0,
       tphlh$SDN$Q = 1.0,
       tphhl$SDN$QN = 1.0,
       tminpwh$CP$D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwl$CP$D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwl$SDN$D_EQ_0 = 1.0,
       tsetup_negedge$D$CP$SDN_EQ_1 = 1.0,
       thold_negedge$D$CP$SDN_EQ_1 = 1.0,
       tsetup_posedge$D$CP$SDN_EQ_1 = 1.0,
       thold_posedge$D$CP$SDN_EQ_1 = 1.0,
       trec$SDN$CP$D_EQ_0 = 1.0,
       trem$SDN$CP$D_EQ_0 = 1.0;

     // path delays
     (posedge CP *> (QN -: D)) = (tpllh$CP$QN, tplhl$CP$QN);
     (posedge CP *> (Q +: D)) = (tpllh$CP$Q, tplhl$CP$Q);
     (negedge SDN *> (QN -: 1'b1)) = (0, tphhl$SDN$QN);
     (negedge SDN *> (Q +: 1'b1)) = (tphlh$SDN$Q, 0);
     $setuphold(posedge CP &&& SDN == 1'b1, negedge D, tsetup_negedge$D$CP$SDN_EQ_1, thold_negedge$D$CP$SDN_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& SDN == 1'b1, posedge D, tsetup_posedge$D$CP$SDN_EQ_1, thold_posedge$D$CP$SDN_EQ_1, NOTIFIER);
     $recrem(posedge SDN, posedge CP &&& D == 1'b0, trec$SDN$CP$D_EQ_0, trem$SDN$CP$D_EQ_0, NOTIFIER);
     $width(posedge CP &&& D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwh$CP$D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(negedge CP &&& D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwl$CP$D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(negedge SDN &&& D == 1'b0, tminpwl$SDN$D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF03HD1 (Q, CP, D, SDN);
input  CP ;
input  D ;
input  SDN ;
output Q ;
reg NOTIFIER ;

   not (I0_SET, SDN);
   udp_dff (N_S_XM21_G, D, CP, 1'B0, I0_SET, NOTIFIER);
   not (N_NET0130_XM18_D, N_S_XM21_G);
   not (Q, N_NET0130_XM18_D);
   not (I5_out, D);
   and (D_EQ_0_AN_SDN_EQ_1, I5_out, SDN);

   specify
     // delay parameters
     specparam
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tphlh$SDN$Q = 1.0,
       tminpwh$CP$D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwl$CP$D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwl$SDN$D_EQ_0 = 1.0,
       tsetup_negedge$D$CP$SDN_EQ_1 = 1.0,
       thold_negedge$D$CP$SDN_EQ_1 = 1.0,
       tsetup_posedge$D$CP$SDN_EQ_1 = 1.0,
       thold_posedge$D$CP$SDN_EQ_1 = 1.0,
       trec$SDN$CP$D_EQ_0 = 1.0,
       trem$SDN$CP$D_EQ_0 = 1.0;

     // path delays
     (posedge CP *> (Q +: D)) = (tpllh$CP$Q, tplhl$CP$Q);
     (negedge SDN *> (Q +: 1'b1)) = (tphlh$SDN$Q, 0);
     $setuphold(posedge CP &&& SDN == 1'b1, negedge D, tsetup_negedge$D$CP$SDN_EQ_1, thold_negedge$D$CP$SDN_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& SDN == 1'b1, posedge D, tsetup_posedge$D$CP$SDN_EQ_1, thold_posedge$D$CP$SDN_EQ_1, NOTIFIER);
     $recrem(posedge SDN, posedge CP &&& D == 1'b0, trec$SDN$CP$D_EQ_0, trem$SDN$CP$D_EQ_0, NOTIFIER);
     $width(posedge CP &&& D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwh$CP$D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(negedge CP &&& D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwl$CP$D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(negedge SDN &&& D == 1'b0, tminpwl$SDN$D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF03HD2 (Q, CP, D, SDN);
input  CP ;
input  D ;
input  SDN ;
output Q ;
reg NOTIFIER ;

   not (I0_SET, SDN);
   udp_dff (N_S_XM21_G, D, CP, 1'B0, I0_SET, NOTIFIER);
   not (N_NET0130_XM18_D, N_S_XM21_G);
   not (Q, N_NET0130_XM18_D);
   not (I5_out, D);
   and (D_EQ_0_AN_SDN_EQ_1, I5_out, SDN);

   specify
     // delay parameters
     specparam
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tphlh$SDN$Q = 1.0,
       tminpwh$CP$D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwl$CP$D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwl$SDN$D_EQ_0 = 1.0,
       tsetup_negedge$D$CP$SDN_EQ_1 = 1.0,
       thold_negedge$D$CP$SDN_EQ_1 = 1.0,
       tsetup_posedge$D$CP$SDN_EQ_1 = 1.0,
       thold_posedge$D$CP$SDN_EQ_1 = 1.0,
       trec$SDN$CP$D_EQ_0 = 1.0,
       trem$SDN$CP$D_EQ_0 = 1.0;

     // path delays
     (posedge CP *> (Q +: D)) = (tpllh$CP$Q, tplhl$CP$Q);
     (negedge SDN *> (Q +: 1'b1)) = (tphlh$SDN$Q, 0);
     $setuphold(posedge CP &&& SDN == 1'b1, negedge D, tsetup_negedge$D$CP$SDN_EQ_1, thold_negedge$D$CP$SDN_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& SDN == 1'b1, posedge D, tsetup_posedge$D$CP$SDN_EQ_1, thold_posedge$D$CP$SDN_EQ_1, NOTIFIER);
     $recrem(posedge SDN, posedge CP &&& D == 1'b0, trec$SDN$CP$D_EQ_0, trem$SDN$CP$D_EQ_0, NOTIFIER);
     $width(posedge CP &&& D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwh$CP$D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(negedge CP &&& D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwl$CP$D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(negedge SDN &&& D == 1'b0, tminpwl$SDN$D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF03HD4 (Q, CP, D, SDN);
input  CP ;
input  D ;
input  SDN ;
output Q ;
reg NOTIFIER ;

   not (I0_SET, SDN);
   udp_dff (N_S_XM21_G, D, CP, 1'B0, I0_SET, NOTIFIER);
   not (N_NET0130_XM18_D, N_S_XM21_G);
   not (Q, N_NET0130_XM18_D);
   not (I5_out, D);
   and (D_EQ_0_AN_SDN_EQ_1, I5_out, SDN);

   specify
     // delay parameters
     specparam
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tphlh$SDN$Q = 1.0,
       tminpwh$CP$D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwl$CP$D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwl$SDN$D_EQ_0 = 1.0,
       tsetup_negedge$D$CP$SDN_EQ_1 = 1.0,
       thold_negedge$D$CP$SDN_EQ_1 = 1.0,
       tsetup_posedge$D$CP$SDN_EQ_1 = 1.0,
       thold_posedge$D$CP$SDN_EQ_1 = 1.0,
       trec$SDN$CP$D_EQ_0 = 1.0,
       trem$SDN$CP$D_EQ_0 = 1.0;

     // path delays
     (posedge CP *> (Q +: D)) = (tpllh$CP$Q, tplhl$CP$Q);
     (negedge SDN *> (Q +: 1'b1)) = (tphlh$SDN$Q, 0);
     $setuphold(posedge CP &&& SDN == 1'b1, negedge D, tsetup_negedge$D$CP$SDN_EQ_1, thold_negedge$D$CP$SDN_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& SDN == 1'b1, posedge D, tsetup_posedge$D$CP$SDN_EQ_1, thold_posedge$D$CP$SDN_EQ_1, NOTIFIER);
     $recrem(posedge SDN, posedge CP &&& D == 1'b0, trec$SDN$CP$D_EQ_0, trem$SDN$CP$D_EQ_0, NOTIFIER);
     $width(posedge CP &&& D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwh$CP$D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(negedge CP &&& D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwl$CP$D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(negedge SDN &&& D == 1'b0, tminpwl$SDN$D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF04D1 (Q, QN, CDN, CP, D, SDN);
input  CDN ;
input  CP ;
input  D ;
input  SDN ;
output Q ;
output QN ;
reg NOTIFIER ;

   not (I0_CLEAR, CDN);
   not (I0_SET, SDN);
   udp_dff (N_S_XM25_G, D, CP, I0_CLEAR, I0_SET, NOTIFIER);
   not (N_NET0130_XM22_D, N_S_XM25_G);
   not (Q, N_NET0130_XM22_D);
   buf (QN, N_NET0130_XM22_D);
   not (I8_out, D);
   and (CDN_EQ_1_AN_D_EQ_0, CDN, I8_out);
   and (CDN_EQ_1_AN_SDN_EQ_1, CDN, SDN);
   and (D_EQ_1_AN_SDN_EQ_1, D, SDN);
   not (I12_out, D);
   and (D_EQ_0_AN_SDN_EQ_1, I12_out, SDN);
   not (I14_out, D);
   and (CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1, CDN, I14_out, SDN);
   not (I17_out, CDN);
   not (I18_out, D);
   and (CDN_EQ_0_AN_D_EQ_0, I17_out, I18_out);

   specify
     // delay parameters
     specparam
       tphhl$CDN$Q = 1.0,
       tphlh$CDN$QN = 1.0,
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tpllh$CP$QN = 1.0,
       tplhl$CP$QN = 1.0,
       tplhl$SDN$Q = 1.0,
       tphlh$SDN$Q = 1.0,
       tpllh$SDN$QN = 1.0,
       tphhl$SDN$QN = 1.0,
       tminpwl$CDN$D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwh$CP$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwl$CP$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwl$SDN$CDN_EQ_0_AN_D_EQ_0 = 1.0,
       tsetup_negedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       thold_negedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       tsetup_posedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       thold_posedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       trec$CDN$CP$D_EQ_1_AN_SDN_EQ_1 = 1.0,
       trem$CDN$CP$D_EQ_1_AN_SDN_EQ_1 = 1.0,
       trec$CDN$SDN$D_EQ_0 = 1.0,
       trec$SDN$CP$CDN_EQ_1_AN_D_EQ_0 = 1.0,
       trem$SDN$CP$CDN_EQ_1_AN_D_EQ_0 = 1.0;

     // path delays
     (posedge CP *> (QN -: D)) = (tpllh$CP$QN, tplhl$CP$QN);
     (posedge CP *> (Q +: D)) = (tpllh$CP$Q, tplhl$CP$Q);
     (negedge SDN *> (QN -: 1'b1)) = (tpllh$SDN$QN, tphhl$SDN$QN);
     (negedge SDN *> (Q +: 1'b1)) = (tphlh$SDN$Q, tplhl$SDN$Q);
     (negedge CDN *> (QN +: 1'b1)) = (tphlh$CDN$QN, 0);
     (negedge CDN *> (Q -: 1'b1)) = (0, tphhl$CDN$Q);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_SDN_EQ_1 == 1'b1, negedge D, tsetup_negedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1, thold_negedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_SDN_EQ_1 == 1'b1, posedge D, tsetup_posedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1, thold_posedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1, NOTIFIER);
     $recrem(posedge CDN, posedge CP &&& D_EQ_1_AN_SDN_EQ_1 == 1'b1, trec$CDN$CP$D_EQ_1_AN_SDN_EQ_1, trem$CDN$CP$D_EQ_1_AN_SDN_EQ_1, NOTIFIER);
     $recovery(posedge CDN, posedge SDN &&& D == 1'b0, trec$CDN$SDN$D_EQ_0, NOTIFIER);
     $recrem(posedge SDN, posedge CP &&& CDN_EQ_1_AN_D_EQ_0 == 1'b1, trec$SDN$CP$CDN_EQ_1_AN_D_EQ_0, trem$SDN$CP$CDN_EQ_1_AN_D_EQ_0, NOTIFIER);
     $width(negedge CDN &&& D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwl$CDN$D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(posedge CP &&& CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwh$CP$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(negedge CP &&& CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwl$CP$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(negedge SDN &&& CDN_EQ_0_AN_D_EQ_0 == 1'b1, tminpwl$SDN$CDN_EQ_0_AN_D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF04D2 (Q, QN, CDN, CP, D, SDN);
input  CDN ;
input  CP ;
input  D ;
input  SDN ;
output Q ;
output QN ;
reg NOTIFIER ;

   not (I0_CLEAR, CDN);
   not (I0_SET, SDN);
   udp_dff (N_S_XM25_G, D, CP, I0_CLEAR, I0_SET, NOTIFIER);
   not (N_NET0130_XM22_D, N_S_XM25_G);
   not (Q, N_NET0130_XM22_D);
   buf (QN, N_NET0130_XM22_D);
   not (I8_out, D);
   and (CDN_EQ_1_AN_D_EQ_0, CDN, I8_out);
   and (CDN_EQ_1_AN_SDN_EQ_1, CDN, SDN);
   and (D_EQ_1_AN_SDN_EQ_1, D, SDN);
   not (I12_out, D);
   and (D_EQ_0_AN_SDN_EQ_1, I12_out, SDN);
   not (I14_out, D);
   and (CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1, CDN, I14_out, SDN);
   not (I17_out, CDN);
   not (I18_out, D);
   and (CDN_EQ_0_AN_D_EQ_0, I17_out, I18_out);

   specify
     // delay parameters
     specparam
       tphhl$CDN$Q = 1.0,
       tphlh$CDN$QN = 1.0,
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tpllh$CP$QN = 1.0,
       tplhl$CP$QN = 1.0,
       tplhl$SDN$Q = 1.0,
       tphlh$SDN$Q = 1.0,
       tpllh$SDN$QN = 1.0,
       tphhl$SDN$QN = 1.0,
       tminpwl$CDN$D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwh$CP$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwl$CP$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwl$SDN$CDN_EQ_0_AN_D_EQ_0 = 1.0,
       tsetup_negedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       thold_negedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       tsetup_posedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       thold_posedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       trec$CDN$CP$D_EQ_1_AN_SDN_EQ_1 = 1.0,
       trem$CDN$CP$D_EQ_1_AN_SDN_EQ_1 = 1.0,
       trec$CDN$SDN$D_EQ_0 = 1.0,
       trec$SDN$CP$CDN_EQ_1_AN_D_EQ_0 = 1.0,
       trem$SDN$CP$CDN_EQ_1_AN_D_EQ_0 = 1.0;

     // path delays
     (posedge CP *> (QN -: D)) = (tpllh$CP$QN, tplhl$CP$QN);
     (posedge CP *> (Q +: D)) = (tpllh$CP$Q, tplhl$CP$Q);
     (negedge SDN *> (QN -: 1'b1)) = (tpllh$SDN$QN, tphhl$SDN$QN);
     (negedge SDN *> (Q +: 1'b1)) = (tphlh$SDN$Q, tplhl$SDN$Q);
     (negedge CDN *> (QN +: 1'b1)) = (tphlh$CDN$QN, 0);
     (negedge CDN *> (Q -: 1'b1)) = (0, tphhl$CDN$Q);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_SDN_EQ_1 == 1'b1, negedge D, tsetup_negedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1, thold_negedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_SDN_EQ_1 == 1'b1, posedge D, tsetup_posedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1, thold_posedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1, NOTIFIER);
     $recrem(posedge CDN, posedge CP &&& D_EQ_1_AN_SDN_EQ_1 == 1'b1, trec$CDN$CP$D_EQ_1_AN_SDN_EQ_1, trem$CDN$CP$D_EQ_1_AN_SDN_EQ_1, NOTIFIER);
     $recovery(posedge CDN, posedge SDN &&& D == 1'b0, trec$CDN$SDN$D_EQ_0, NOTIFIER);
     $recrem(posedge SDN, posedge CP &&& CDN_EQ_1_AN_D_EQ_0 == 1'b1, trec$SDN$CP$CDN_EQ_1_AN_D_EQ_0, trem$SDN$CP$CDN_EQ_1_AN_D_EQ_0, NOTIFIER);
     $width(negedge CDN &&& D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwl$CDN$D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(posedge CP &&& CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwh$CP$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(negedge CP &&& CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwl$CP$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(negedge SDN &&& CDN_EQ_0_AN_D_EQ_0 == 1'b1, tminpwl$SDN$CDN_EQ_0_AN_D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF04D4 (Q, QN, CDN, CP, D, SDN);
input  CDN ;
input  CP ;
input  D ;
input  SDN ;
output Q ;
output QN ;
reg NOTIFIER ;

   not (I0_CLEAR, CDN);
   not (I0_SET, SDN);
   udp_dff (N_S_XM25_G, D, CP, I0_CLEAR, I0_SET, NOTIFIER);
   not (N_NET0130_XM22_D, N_S_XM25_G);
   not (Q, N_NET0130_XM22_D);
   buf (QN, N_NET0130_XM22_D);
   not (I8_out, D);
   and (CDN_EQ_1_AN_D_EQ_0, CDN, I8_out);
   and (CDN_EQ_1_AN_SDN_EQ_1, CDN, SDN);
   and (D_EQ_1_AN_SDN_EQ_1, D, SDN);
   not (I12_out, D);
   and (D_EQ_0_AN_SDN_EQ_1, I12_out, SDN);
   not (I14_out, D);
   and (CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1, CDN, I14_out, SDN);
   not (I17_out, CDN);
   not (I18_out, D);
   and (CDN_EQ_0_AN_D_EQ_0, I17_out, I18_out);

   specify
     // delay parameters
     specparam
       tphhl$CDN$Q = 1.0,
       tphlh$CDN$QN = 1.0,
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tpllh$CP$QN = 1.0,
       tplhl$CP$QN = 1.0,
       tplhl$SDN$Q = 1.0,
       tphlh$SDN$Q = 1.0,
       tpllh$SDN$QN = 1.0,
       tphhl$SDN$QN = 1.0,
       tminpwl$CDN$D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwh$CP$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwl$CP$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwl$SDN$CDN_EQ_0_AN_D_EQ_0 = 1.0,
       tsetup_negedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       thold_negedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       tsetup_posedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       thold_posedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       trec$CDN$CP$D_EQ_1_AN_SDN_EQ_1 = 1.0,
       trem$CDN$CP$D_EQ_1_AN_SDN_EQ_1 = 1.0,
       trec$CDN$SDN$D_EQ_0 = 1.0,
       trec$SDN$CP$CDN_EQ_1_AN_D_EQ_0 = 1.0,
       trem$SDN$CP$CDN_EQ_1_AN_D_EQ_0 = 1.0;

     // path delays
     (posedge CP *> (QN -: D)) = (tpllh$CP$QN, tplhl$CP$QN);
     (posedge CP *> (Q +: D)) = (tpllh$CP$Q, tplhl$CP$Q);
     (negedge SDN *> (QN -: 1'b1)) = (tpllh$SDN$QN, tphhl$SDN$QN);
     (negedge SDN *> (Q +: 1'b1)) = (tphlh$SDN$Q, tplhl$SDN$Q);
     (negedge CDN *> (QN +: 1'b1)) = (tphlh$CDN$QN, 0);
     (negedge CDN *> (Q -: 1'b1)) = (0, tphhl$CDN$Q);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_SDN_EQ_1 == 1'b1, negedge D, tsetup_negedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1, thold_negedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_SDN_EQ_1 == 1'b1, posedge D, tsetup_posedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1, thold_posedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1, NOTIFIER);
     $recrem(posedge CDN, posedge CP &&& D_EQ_1_AN_SDN_EQ_1 == 1'b1, trec$CDN$CP$D_EQ_1_AN_SDN_EQ_1, trem$CDN$CP$D_EQ_1_AN_SDN_EQ_1, NOTIFIER);
     $recovery(posedge CDN, posedge SDN &&& D == 1'b0, trec$CDN$SDN$D_EQ_0, NOTIFIER);
     $recrem(posedge SDN, posedge CP &&& CDN_EQ_1_AN_D_EQ_0 == 1'b1, trec$SDN$CP$CDN_EQ_1_AN_D_EQ_0, trem$SDN$CP$CDN_EQ_1_AN_D_EQ_0, NOTIFIER);
     $width(negedge CDN &&& D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwl$CDN$D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(posedge CP &&& CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwh$CP$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(negedge CP &&& CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwl$CP$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(negedge SDN &&& CDN_EQ_0_AN_D_EQ_0 == 1'b1, tminpwl$SDN$CDN_EQ_0_AN_D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF05D1 (Q, QN, CPN, D);
input  CPN ;
input  D ;
output Q ;
output QN ;
reg NOTIFIER ;
reg ReSeT;
`ifdef  RSTn_lib
   
	 initial begin
		ReSeT = 0 ;
		#3 ReSeT = 1 ;
		#111 ReSeT = 0 ;
	end
  `else initial  ReSeT = 0;
`endif
   not (I0_CLOCK, CPN);
   udp_dff (N_S_XM19_G, D, I0_CLOCK, ReSeT , 1'B0, NOTIFIER);

   not (N_NET0130_XM16_D, N_S_XM19_G);
   buf (Q, N_S_XM19_G);
   not (QN, N_S_XM19_G);

   specify
     // delay parameters
     specparam
       tphlh$CPN$Q = 1.0,
       tphhl$CPN$Q = 1.0,
       tphlh$CPN$QN = 1.0,
       tphhl$CPN$QN = 1.0,
       tminpwh$CPN$D_EQ_0 = 1.0,
       tminpwl$CPN$D_EQ_0 = 1.0,
       tsetup_negedge$D$CPN = 1.0,
       thold_negedge$D$CPN = 1.0,
       tsetup_posedge$D$CPN = 1.0,
       thold_posedge$D$CPN = 1.0;

     // path delays
     (negedge CPN *> (QN -: D)) = (tphlh$CPN$QN, tphhl$CPN$QN);
     (negedge CPN *> (Q +: D)) = (tphlh$CPN$Q, tphhl$CPN$Q);
     $setuphold(negedge CPN, negedge D, tsetup_negedge$D$CPN, thold_negedge$D$CPN, NOTIFIER);
     $setuphold(negedge CPN, posedge D, tsetup_posedge$D$CPN, thold_posedge$D$CPN, NOTIFIER);
     $width(posedge CPN &&& D == 1'b0, tminpwh$CPN$D_EQ_0, 0, NOTIFIER);
     $width(negedge CPN &&& D == 1'b0, tminpwl$CPN$D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF05D2 (Q, QN, CPN, D);
input  CPN ;
input  D ;
output Q ;
output QN ;
reg NOTIFIER ;

   not (I0_CLOCK, CPN);
   udp_dff (N_S_XM19_G, D, I0_CLOCK, 1'B0, 1'B0, NOTIFIER);
   not (N_NET0130_XM16_D, N_S_XM19_G);
   buf (Q, N_S_XM19_G);
   not (QN, N_S_XM19_G);

   specify
     // delay parameters
     specparam
       tphlh$CPN$Q = 1.0,
       tphhl$CPN$Q = 1.0,
       tphlh$CPN$QN = 1.0,
       tphhl$CPN$QN = 1.0,
       tminpwh$CPN$D_EQ_0 = 1.0,
       tminpwl$CPN$D_EQ_0 = 1.0,
       tsetup_negedge$D$CPN = 1.0,
       thold_negedge$D$CPN = 1.0,
       tsetup_posedge$D$CPN = 1.0,
       thold_posedge$D$CPN = 1.0;

     // path delays
     (negedge CPN *> (QN -: D)) = (tphlh$CPN$QN, tphhl$CPN$QN);
     (negedge CPN *> (Q +: D)) = (tphlh$CPN$Q, tphhl$CPN$Q);
     $setuphold(negedge CPN, negedge D, tsetup_negedge$D$CPN, thold_negedge$D$CPN, NOTIFIER);
     $setuphold(negedge CPN, posedge D, tsetup_posedge$D$CPN, thold_posedge$D$CPN, NOTIFIER);
     $width(posedge CPN &&& D == 1'b0, tminpwh$CPN$D_EQ_0, 0, NOTIFIER);
     $width(negedge CPN &&& D == 1'b0, tminpwl$CPN$D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF05D4 (Q, QN, CPN, D);
input  CPN ;
input  D ;
output Q ;
output QN ;
reg NOTIFIER ;

   not (I0_CLOCK, CPN);
   udp_dff (N_S_XM19_G, D, I0_CLOCK, 1'B0, 1'B0, NOTIFIER);
   not (N_NET0130_XM16_D, N_S_XM19_G);
   buf (Q, N_S_XM19_G);
   not (QN, N_S_XM19_G);

   specify
     // delay parameters
     specparam
       tphlh$CPN$Q = 1.0,
       tphhl$CPN$Q = 1.0,
       tphlh$CPN$QN = 1.0,
       tphhl$CPN$QN = 1.0,
       tminpwh$CPN$D_EQ_0 = 1.0,
       tminpwl$CPN$D_EQ_0 = 1.0,
       tsetup_negedge$D$CPN = 1.0,
       thold_negedge$D$CPN = 1.0,
       tsetup_posedge$D$CPN = 1.0,
       thold_posedge$D$CPN = 1.0;

     // path delays
     (negedge CPN *> (QN -: D)) = (tphlh$CPN$QN, tphhl$CPN$QN);
     (negedge CPN *> (Q +: D)) = (tphlh$CPN$Q, tphhl$CPN$Q);
     $setuphold(negedge CPN, negedge D, tsetup_negedge$D$CPN, thold_negedge$D$CPN, NOTIFIER);
     $setuphold(negedge CPN, posedge D, tsetup_posedge$D$CPN, thold_posedge$D$CPN, NOTIFIER);
     $width(posedge CPN &&& D == 1'b0, tminpwh$CPN$D_EQ_0, 0, NOTIFIER);
     $width(negedge CPN &&& D == 1'b0, tminpwl$CPN$D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF05ED1 (Q, QN, CPN, D, E);
input  CPN ;
input  D ;
input  E ;
output Q ;
output QN ;
reg NOTIFIER ;

   udp_mux2 (I0_D, N_S_XM3_G, D, E);
   not (I0_CLOCK, CPN);
   udp_dff (N_S_XM3_G, I0_D, I0_CLOCK, 1'B0, 1'B0, NOTIFIER);
   not (N_NET0235_XM29_G, N_S_XM3_G);
   not (Q, N_NET0235_XM29_G);
   buf (QN, N_NET0235_XM29_G);
   not (I8_out, D);
   and (D_EQ_0_AN_E_EQ_1, I8_out, E);

   specify
     // delay parameters
     specparam
       tphlh$CPN$Q = 1.0,
       tphhl$CPN$Q = 1.0,
       tphlh$CPN$QN = 1.0,
       tphhl$CPN$QN = 1.0,
       tminpwh$CPN$D_EQ_0_AN_E_EQ_1 = 1.0,
       tminpwl$CPN$D_EQ_0_AN_E_EQ_1 = 1.0,
       tsetup_negedge$D$CPN$E_EQ_1 = 1.0,
       thold_negedge$D$CPN$E_EQ_1 = 1.0,
       tsetup_negedge$E$CPN$D_EQ_0 = 1.0,
       thold_negedge$E$CPN$D_EQ_0 = 1.0,
       tsetup_negedge$E$CPN$D_EQ_1 = 1.0,
       thold_negedge$E$CPN$D_EQ_1 = 1.0,
       tsetup_posedge$D$CPN$E_EQ_1 = 1.0,
       thold_posedge$D$CPN$E_EQ_1 = 1.0,
       tsetup_posedge$E$CPN$D_EQ_0 = 1.0,
       thold_posedge$E$CPN$D_EQ_0 = 1.0,
       tsetup_posedge$E$CPN$D_EQ_1 = 1.0,
       thold_posedge$E$CPN$D_EQ_1 = 1.0;

     // path delays
     (negedge CPN *> (QN -: E?D:N_S_XM3_G)) = (tphlh$CPN$QN, tphhl$CPN$QN);
     (negedge CPN *> (Q +: E?D:N_S_XM3_G)) = (tphlh$CPN$Q, tphhl$CPN$Q);
     $setuphold(negedge CPN &&& E == 1'b1, negedge D, tsetup_negedge$D$CPN$E_EQ_1, thold_negedge$D$CPN$E_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& D == 1'b0, negedge E, tsetup_negedge$E$CPN$D_EQ_0, thold_negedge$E$CPN$D_EQ_0, NOTIFIER);
     $setuphold(negedge CPN &&& D == 1'b1, negedge E, tsetup_negedge$E$CPN$D_EQ_1, thold_negedge$E$CPN$D_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& E == 1'b1, posedge D, tsetup_posedge$D$CPN$E_EQ_1, thold_posedge$D$CPN$E_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& D == 1'b0, posedge E, tsetup_posedge$E$CPN$D_EQ_0, thold_posedge$E$CPN$D_EQ_0, NOTIFIER);
     $setuphold(negedge CPN &&& D == 1'b1, posedge E, tsetup_posedge$E$CPN$D_EQ_1, thold_posedge$E$CPN$D_EQ_1, NOTIFIER);
     $width(posedge CPN &&& D_EQ_0_AN_E_EQ_1 == 1'b1, tminpwh$CPN$D_EQ_0_AN_E_EQ_1, 0, NOTIFIER);
     $width(negedge CPN &&& D_EQ_0_AN_E_EQ_1 == 1'b1, tminpwl$CPN$D_EQ_0_AN_E_EQ_1, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF05ED2 (Q, QN, CPN, D, E);
input  CPN ;
input  D ;
input  E ;
output Q ;
output QN ;
reg NOTIFIER ;

   udp_mux2 (I0_D, N_S_XM3_G, D, E);
   not (I0_CLOCK, CPN);
   udp_dff (N_S_XM3_G, I0_D, I0_CLOCK, 1'B0, 1'B0, NOTIFIER);
   not (N_NET0235_XM29_G, N_S_XM3_G);
   not (Q, N_NET0235_XM29_G);
   buf (QN, N_NET0235_XM29_G);
   not (I8_out, D);
   and (D_EQ_0_AN_E_EQ_1, I8_out, E);

   specify
     // delay parameters
     specparam
       tphlh$CPN$Q = 1.0,
       tphhl$CPN$Q = 1.0,
       tphlh$CPN$QN = 1.0,
       tphhl$CPN$QN = 1.0,
       tminpwh$CPN$D_EQ_0_AN_E_EQ_1 = 1.0,
       tminpwl$CPN$D_EQ_0_AN_E_EQ_1 = 1.0,
       tsetup_negedge$D$CPN$E_EQ_1 = 1.0,
       thold_negedge$D$CPN$E_EQ_1 = 1.0,
       tsetup_negedge$E$CPN$D_EQ_0 = 1.0,
       thold_negedge$E$CPN$D_EQ_0 = 1.0,
       tsetup_negedge$E$CPN$D_EQ_1 = 1.0,
       thold_negedge$E$CPN$D_EQ_1 = 1.0,
       tsetup_posedge$D$CPN$E_EQ_1 = 1.0,
       thold_posedge$D$CPN$E_EQ_1 = 1.0,
       tsetup_posedge$E$CPN$D_EQ_0 = 1.0,
       thold_posedge$E$CPN$D_EQ_0 = 1.0,
       tsetup_posedge$E$CPN$D_EQ_1 = 1.0,
       thold_posedge$E$CPN$D_EQ_1 = 1.0;

     // path delays
     (negedge CPN *> (QN -: E?D:N_S_XM3_G)) = (tphlh$CPN$QN, tphhl$CPN$QN);
     (negedge CPN *> (Q +: E?D:N_S_XM3_G)) = (tphlh$CPN$Q, tphhl$CPN$Q);
     $setuphold(negedge CPN &&& E == 1'b1, negedge D, tsetup_negedge$D$CPN$E_EQ_1, thold_negedge$D$CPN$E_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& D == 1'b0, negedge E, tsetup_negedge$E$CPN$D_EQ_0, thold_negedge$E$CPN$D_EQ_0, NOTIFIER);
     $setuphold(negedge CPN &&& D == 1'b1, negedge E, tsetup_negedge$E$CPN$D_EQ_1, thold_negedge$E$CPN$D_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& E == 1'b1, posedge D, tsetup_posedge$D$CPN$E_EQ_1, thold_posedge$D$CPN$E_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& D == 1'b0, posedge E, tsetup_posedge$E$CPN$D_EQ_0, thold_posedge$E$CPN$D_EQ_0, NOTIFIER);
     $setuphold(negedge CPN &&& D == 1'b1, posedge E, tsetup_posedge$E$CPN$D_EQ_1, thold_posedge$E$CPN$D_EQ_1, NOTIFIER);
     $width(posedge CPN &&& D_EQ_0_AN_E_EQ_1 == 1'b1, tminpwh$CPN$D_EQ_0_AN_E_EQ_1, 0, NOTIFIER);
     $width(negedge CPN &&& D_EQ_0_AN_E_EQ_1 == 1'b1, tminpwl$CPN$D_EQ_0_AN_E_EQ_1, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF05ED4 (Q, QN, CPN, D, E);
input  CPN ;
input  D ;
input  E ;
output Q ;
output QN ;
reg NOTIFIER ;

   udp_mux2 (I0_D, N_S_XM3_G, D, E);
   not (I0_CLOCK, CPN);
   udp_dff (N_S_XM3_G, I0_D, I0_CLOCK, 1'B0, 1'B0, NOTIFIER);
   not (N_NET0235_XM29_G, N_S_XM3_G);
   not (Q, N_NET0235_XM29_G);
   buf (QN, N_NET0235_XM29_G);
   not (I8_out, D);
   and (D_EQ_0_AN_E_EQ_1, I8_out, E);

   specify
     // delay parameters
     specparam
       tphlh$CPN$Q = 1.0,
       tphhl$CPN$Q = 1.0,
       tphlh$CPN$QN = 1.0,
       tphhl$CPN$QN = 1.0,
       tminpwh$CPN$D_EQ_0_AN_E_EQ_1 = 1.0,
       tminpwl$CPN$D_EQ_0_AN_E_EQ_1 = 1.0,
       tsetup_negedge$D$CPN$E_EQ_1 = 1.0,
       thold_negedge$D$CPN$E_EQ_1 = 1.0,
       tsetup_negedge$E$CPN$D_EQ_0 = 1.0,
       thold_negedge$E$CPN$D_EQ_0 = 1.0,
       tsetup_negedge$E$CPN$D_EQ_1 = 1.0,
       thold_negedge$E$CPN$D_EQ_1 = 1.0,
       tsetup_posedge$D$CPN$E_EQ_1 = 1.0,
       thold_posedge$D$CPN$E_EQ_1 = 1.0,
       tsetup_posedge$E$CPN$D_EQ_0 = 1.0,
       thold_posedge$E$CPN$D_EQ_0 = 1.0,
       tsetup_posedge$E$CPN$D_EQ_1 = 1.0,
       thold_posedge$E$CPN$D_EQ_1 = 1.0;

     // path delays
     (negedge CPN *> (QN -: E?D:N_S_XM3_G)) = (tphlh$CPN$QN, tphhl$CPN$QN);
     (negedge CPN *> (Q +: E?D:N_S_XM3_G)) = (tphlh$CPN$Q, tphhl$CPN$Q);
     $setuphold(negedge CPN &&& E == 1'b1, negedge D, tsetup_negedge$D$CPN$E_EQ_1, thold_negedge$D$CPN$E_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& D == 1'b0, negedge E, tsetup_negedge$E$CPN$D_EQ_0, thold_negedge$E$CPN$D_EQ_0, NOTIFIER);
     $setuphold(negedge CPN &&& D == 1'b1, negedge E, tsetup_negedge$E$CPN$D_EQ_1, thold_negedge$E$CPN$D_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& E == 1'b1, posedge D, tsetup_posedge$D$CPN$E_EQ_1, thold_posedge$D$CPN$E_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& D == 1'b0, posedge E, tsetup_posedge$E$CPN$D_EQ_0, thold_posedge$E$CPN$D_EQ_0, NOTIFIER);
     $setuphold(negedge CPN &&& D == 1'b1, posedge E, tsetup_posedge$E$CPN$D_EQ_1, thold_posedge$E$CPN$D_EQ_1, NOTIFIER);
     $width(posedge CPN &&& D_EQ_0_AN_E_EQ_1 == 1'b1, tminpwh$CPN$D_EQ_0_AN_E_EQ_1, 0, NOTIFIER);
     $width(negedge CPN &&& D_EQ_0_AN_E_EQ_1 == 1'b1, tminpwl$CPN$D_EQ_0_AN_E_EQ_1, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF05HD1 (Q, CPN, D);
input  CPN ;
input  D ;
output Q ;
reg NOTIFIER ;
reg ReSeT;

 `ifdef  RSTn_lib
    
	 initial begin
		ReSeT = 0 ;
		#3 ReSeT = 1 ;
		#111 ReSeT = 0 ;
	end

  `else initial  ReSeT = 0;
`endif
   not (I0_CLOCK, CPN);
   udp_dff (N_S_XM19_G, D, I0_CLOCK, ReSeT, 1'B0, NOTIFIER);
   not (N_NET0130_XM16_D, N_S_XM19_G);
   buf (Q, N_S_XM19_G);

   specify
     // delay parameters
     specparam
       tphlh$CPN$Q = 1.0,
       tphhl$CPN$Q = 1.0,
       tminpwh$CPN$D_EQ_0 = 1.0,
       tminpwl$CPN$D_EQ_0 = 1.0,
       tsetup_negedge$D$CPN = 1.0,
       thold_negedge$D$CPN = 1.0,
       tsetup_posedge$D$CPN = 1.0,
       thold_posedge$D$CPN = 1.0;

     // path delays
     (negedge CPN *> (Q +: D)) = (tphlh$CPN$Q, tphhl$CPN$Q);
     $setuphold(negedge CPN, negedge D, tsetup_negedge$D$CPN, thold_negedge$D$CPN, NOTIFIER);
     $setuphold(negedge CPN, posedge D, tsetup_posedge$D$CPN, thold_posedge$D$CPN, NOTIFIER);
     $width(posedge CPN &&& D == 1'b0, tminpwh$CPN$D_EQ_0, 0, NOTIFIER);
     $width(negedge CPN &&& D == 1'b0, tminpwl$CPN$D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF05HD2 (Q, CPN, D);
input  CPN ;
input  D ;
output Q ;
reg NOTIFIER ;
reg ReSeT;
 
`ifdef  RSTn_lib
	 initial begin
		ReSeT = 0 ;
		#3 ReSeT = 1 ;
		#111 ReSeT = 0 ;
	end
  `else initial  ReSeT = 0;
`endif
   not (I0_CLOCK, CPN);
   udp_dff (N_S_XM19_G, D, I0_CLOCK, ReSeT, 1'B0, NOTIFIER);

   not (N_NET0130_XM16_D, N_S_XM19_G);
   buf (Q, N_S_XM19_G);

   specify
     // delay parameters
     specparam
       tphlh$CPN$Q = 1.0,
       tphhl$CPN$Q = 1.0,
       tminpwh$CPN$D_EQ_0 = 1.0,
       tminpwl$CPN$D_EQ_0 = 1.0,
       tsetup_negedge$D$CPN = 1.0,
       thold_negedge$D$CPN = 1.0,
       tsetup_posedge$D$CPN = 1.0,
       thold_posedge$D$CPN = 1.0;

     // path delays
     (negedge CPN *> (Q +: D)) = (tphlh$CPN$Q, tphhl$CPN$Q);
     $setuphold(negedge CPN, negedge D, tsetup_negedge$D$CPN, thold_negedge$D$CPN, NOTIFIER);
     $setuphold(negedge CPN, posedge D, tsetup_posedge$D$CPN, thold_posedge$D$CPN, NOTIFIER);
     $width(posedge CPN &&& D == 1'b0, tminpwh$CPN$D_EQ_0, 0, NOTIFIER);
     $width(negedge CPN &&& D == 1'b0, tminpwl$CPN$D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF05HD4 (Q, CPN, D);
input  CPN ;
input  D ;
output Q ;
reg NOTIFIER ;
reg ReSeT;

 `ifdef  RSTn_lib
	 initial begin
		ReSeT = 0 ;
		#3 ReSeT = 1 ;
		#111 ReSeT = 0 ;
	end
  `else initial  ReSeT = 0;
`endif

   not (I0_CLOCK, CPN);
   udp_dff (N_S_XM19_G, D, I0_CLOCK, ReSeT, 1'B0, NOTIFIER);

   not (N_NET0130_XM16_D, N_S_XM19_G);
   buf (Q, N_S_XM19_G);

   specify
     // delay parameters
     specparam
       tphlh$CPN$Q = 1.0,
       tphhl$CPN$Q = 1.0,
       tminpwh$CPN$D_EQ_0 = 1.0,
       tminpwl$CPN$D_EQ_0 = 1.0,
       tsetup_negedge$D$CPN = 1.0,
       thold_negedge$D$CPN = 1.0,
       tsetup_posedge$D$CPN = 1.0,
       thold_posedge$D$CPN = 1.0;

     // path delays
     (negedge CPN *> (Q +: D)) = (tphlh$CPN$Q, tphhl$CPN$Q);
     $setuphold(negedge CPN, negedge D, tsetup_negedge$D$CPN, thold_negedge$D$CPN, NOTIFIER);
     $setuphold(negedge CPN, posedge D, tsetup_posedge$D$CPN, thold_posedge$D$CPN, NOTIFIER);
     $width(posedge CPN &&& D == 1'b0, tminpwh$CPN$D_EQ_0, 0, NOTIFIER);
     $width(negedge CPN &&& D == 1'b0, tminpwl$CPN$D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF06D1 (Q, QN, CDN, CPN, D);
input  CDN ;
input  CPN ;
input  D ;
output Q ;
output QN ;
reg NOTIFIER ;

   not (I0_CLOCK, CPN);
   not (I0_CLEAR, CDN);
   udp_dff (N_S_XM23_G, D, I0_CLOCK, I0_CLEAR, 1'B0, NOTIFIER);
   not (N_NET0130_XM20_D, N_S_XM23_G);
   buf (Q, N_S_XM23_G);
   not (QN, N_S_XM23_G);
   not (I8_out, D);
   and (CDN_EQ_1_AN_D_EQ_0, CDN, I8_out);

   specify
     // delay parameters
     specparam
       tphhl$CDN$Q = 1.0,
       tphlh$CDN$QN = 1.0,
       tphlh$CPN$Q = 1.0,
       tphhl$CPN$Q = 1.0,
       tphlh$CPN$QN = 1.0,
       tphhl$CPN$QN = 1.0,
       tminpwl$CDN$D_EQ_0 = 1.0,
       tminpwh$CPN$CDN_EQ_1_AN_D_EQ_0 = 1.0,
       tminpwl$CPN$CDN_EQ_1_AN_D_EQ_0 = 1.0,
       tsetup_negedge$D$CPN$CDN_EQ_1 = 1.0,
       thold_negedge$D$CPN$CDN_EQ_1 = 1.0,
       tsetup_posedge$D$CPN$CDN_EQ_1 = 1.0,
       thold_posedge$D$CPN$CDN_EQ_1 = 1.0,
       trec$CDN$CPN$D_EQ_1 = 1.0,
       trem$CDN$CPN$D_EQ_1 = 1.0;

     // path delays
     (negedge CPN *> (QN -: D)) = (tphlh$CPN$QN, tphhl$CPN$QN);
     (negedge CPN *> (Q +: D)) = (tphlh$CPN$Q, tphhl$CPN$Q);
     (negedge CDN *> (QN +: 1'b1)) = (tphlh$CDN$QN, 0);
     (negedge CDN *> (Q -: 1'b1)) = (0, tphhl$CDN$Q);
     $setuphold(negedge CPN &&& CDN == 1'b1, negedge D, tsetup_negedge$D$CPN$CDN_EQ_1, thold_negedge$D$CPN$CDN_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& CDN == 1'b1, posedge D, tsetup_posedge$D$CPN$CDN_EQ_1, thold_posedge$D$CPN$CDN_EQ_1, NOTIFIER);
     $recrem(posedge CDN, negedge CPN &&& D == 1'b1, trec$CDN$CPN$D_EQ_1, trem$CDN$CPN$D_EQ_1, NOTIFIER);
     $width(negedge CDN &&& D == 1'b0, tminpwl$CDN$D_EQ_0, 0, NOTIFIER);
     $width(posedge CPN &&& CDN_EQ_1_AN_D_EQ_0 == 1'b1, tminpwh$CPN$CDN_EQ_1_AN_D_EQ_0, 0, NOTIFIER);
     $width(negedge CPN &&& CDN_EQ_1_AN_D_EQ_0 == 1'b1, tminpwl$CPN$CDN_EQ_1_AN_D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF06D2 (Q, QN, CDN, CPN, D);
input  CDN ;
input  CPN ;
input  D ;
output Q ;
output QN ;
reg NOTIFIER ;

   not (I0_CLOCK, CPN);
   not (I0_CLEAR, CDN);
   udp_dff (N_S_XM23_G, D, I0_CLOCK, I0_CLEAR, 1'B0, NOTIFIER);
   not (N_NET0130_XM20_D, N_S_XM23_G);
   buf (Q, N_S_XM23_G);
   not (QN, N_S_XM23_G);
   not (I8_out, D);
   and (CDN_EQ_1_AN_D_EQ_0, CDN, I8_out);

   specify
     // delay parameters
     specparam
       tphhl$CDN$Q = 1.0,
       tphlh$CDN$QN = 1.0,
       tphlh$CPN$Q = 1.0,
       tphhl$CPN$Q = 1.0,
       tphlh$CPN$QN = 1.0,
       tphhl$CPN$QN = 1.0,
       tminpwl$CDN$D_EQ_0 = 1.0,
       tminpwh$CPN$CDN_EQ_1_AN_D_EQ_0 = 1.0,
       tminpwl$CPN$CDN_EQ_1_AN_D_EQ_0 = 1.0,
       tsetup_negedge$D$CPN$CDN_EQ_1 = 1.0,
       thold_negedge$D$CPN$CDN_EQ_1 = 1.0,
       tsetup_posedge$D$CPN$CDN_EQ_1 = 1.0,
       thold_posedge$D$CPN$CDN_EQ_1 = 1.0,
       trec$CDN$CPN$D_EQ_1 = 1.0,
       trem$CDN$CPN$D_EQ_1 = 1.0;

     // path delays
     (negedge CPN *> (QN -: D)) = (tphlh$CPN$QN, tphhl$CPN$QN);
     (negedge CPN *> (Q +: D)) = (tphlh$CPN$Q, tphhl$CPN$Q);
     (negedge CDN *> (QN +: 1'b1)) = (tphlh$CDN$QN, 0);
     (negedge CDN *> (Q -: 1'b1)) = (0, tphhl$CDN$Q);
     $setuphold(negedge CPN &&& CDN == 1'b1, negedge D, tsetup_negedge$D$CPN$CDN_EQ_1, thold_negedge$D$CPN$CDN_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& CDN == 1'b1, posedge D, tsetup_posedge$D$CPN$CDN_EQ_1, thold_posedge$D$CPN$CDN_EQ_1, NOTIFIER);
     $recrem(posedge CDN, negedge CPN &&& D == 1'b1, trec$CDN$CPN$D_EQ_1, trem$CDN$CPN$D_EQ_1, NOTIFIER);
     $width(negedge CDN &&& D == 1'b0, tminpwl$CDN$D_EQ_0, 0, NOTIFIER);
     $width(posedge CPN &&& CDN_EQ_1_AN_D_EQ_0 == 1'b1, tminpwh$CPN$CDN_EQ_1_AN_D_EQ_0, 0, NOTIFIER);
     $width(negedge CPN &&& CDN_EQ_1_AN_D_EQ_0 == 1'b1, tminpwl$CPN$CDN_EQ_1_AN_D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF06D4 (Q, QN, CDN, CPN, D);
input  CDN ;
input  CPN ;
input  D ;
output Q ;
output QN ;
reg NOTIFIER ;

   not (I0_CLOCK, CPN);
   not (I0_CLEAR, CDN);
   udp_dff (N_S_XM23_G, D, I0_CLOCK, I0_CLEAR, 1'B0, NOTIFIER);
   not (N_NET0130_XM20_D, N_S_XM23_G);
   buf (Q, N_S_XM23_G);
   not (QN, N_S_XM23_G);
   not (I8_out, D);
   and (CDN_EQ_1_AN_D_EQ_0, CDN, I8_out);

   specify
     // delay parameters
     specparam
       tphhl$CDN$Q = 1.0,
       tphlh$CDN$QN = 1.0,
       tphlh$CPN$Q = 1.0,
       tphhl$CPN$Q = 1.0,
       tphlh$CPN$QN = 1.0,
       tphhl$CPN$QN = 1.0,
       tminpwl$CDN$D_EQ_0 = 1.0,
       tminpwh$CPN$CDN_EQ_1_AN_D_EQ_0 = 1.0,
       tminpwl$CPN$CDN_EQ_1_AN_D_EQ_0 = 1.0,
       tsetup_negedge$D$CPN$CDN_EQ_1 = 1.0,
       thold_negedge$D$CPN$CDN_EQ_1 = 1.0,
       tsetup_posedge$D$CPN$CDN_EQ_1 = 1.0,
       thold_posedge$D$CPN$CDN_EQ_1 = 1.0,
       trec$CDN$CPN$D_EQ_1 = 1.0,
       trem$CDN$CPN$D_EQ_1 = 1.0;

     // path delays
     (negedge CPN *> (QN -: D)) = (tphlh$CPN$QN, tphhl$CPN$QN);
     (negedge CPN *> (Q +: D)) = (tphlh$CPN$Q, tphhl$CPN$Q);
     (negedge CDN *> (QN +: 1'b1)) = (tphlh$CDN$QN, 0);
     (negedge CDN *> (Q -: 1'b1)) = (0, tphhl$CDN$Q);
     $setuphold(negedge CPN &&& CDN == 1'b1, negedge D, tsetup_negedge$D$CPN$CDN_EQ_1, thold_negedge$D$CPN$CDN_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& CDN == 1'b1, posedge D, tsetup_posedge$D$CPN$CDN_EQ_1, thold_posedge$D$CPN$CDN_EQ_1, NOTIFIER);
     $recrem(posedge CDN, negedge CPN &&& D == 1'b1, trec$CDN$CPN$D_EQ_1, trem$CDN$CPN$D_EQ_1, NOTIFIER);
     $width(negedge CDN &&& D == 1'b0, tminpwl$CDN$D_EQ_0, 0, NOTIFIER);
     $width(posedge CPN &&& CDN_EQ_1_AN_D_EQ_0 == 1'b1, tminpwh$CPN$CDN_EQ_1_AN_D_EQ_0, 0, NOTIFIER);
     $width(negedge CPN &&& CDN_EQ_1_AN_D_EQ_0 == 1'b1, tminpwl$CPN$CDN_EQ_1_AN_D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF06ED1 (Q, QN, CDN, CPN, D, E);
input  CDN ;
input  CPN ;
input  D ;
input  E ;
output Q ;
output QN ;
reg NOTIFIER ;

   udp_mux2 (I0_D, N_S_XM3_G, D, E);
   not (I0_CLOCK, CPN);
   not (I0_CLEAR, CDN);
   udp_dff (N_S_XM3_G, I0_D, I0_CLOCK, I0_CLEAR, 1'B0, NOTIFIER);
   not (N_NET0235_XM31_G, N_S_XM3_G);
   not (Q, N_NET0235_XM31_G);
   not (QN, N_S_XM3_G);
   and (CDN_EQ_1_AN_E_EQ_1, CDN, E);
   and (D_EQ_1_AN_E_EQ_1, D, E);
   not (I10_out, D);
   not (I11_out, E);
   and (D_EQ_0_AN_E_EQ_0, I10_out, I11_out);
   not (I13_out, D);
   and (CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1, CDN, I13_out, E);

   specify
     // delay parameters
     specparam
       tphhl$CDN$Q = 1.0,
       tphlh$CDN$QN = 1.0,
       tphlh$CPN$Q = 1.0,
       tphhl$CPN$Q = 1.0,
       tphlh$CPN$QN = 1.0,
       tphhl$CPN$QN = 1.0,
       tminpwl$CDN$D_EQ_0_AN_E_EQ_0 = 1.0,
       tminpwh$CPN$CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1 = 1.0,
       tminpwl$CPN$CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1 = 1.0,
       tsetup_negedge$D$CPN$CDN_EQ_1_AN_E_EQ_1 = 1.0,
       thold_negedge$D$CPN$CDN_EQ_1_AN_E_EQ_1 = 1.0,
       tsetup_negedge$E$CPN$CDN_EQ_1 = 1.0,
       thold_negedge$E$CPN$CDN_EQ_1 = 1.0,
       tsetup_posedge$D$CPN$CDN_EQ_1_AN_E_EQ_1 = 1.0,
       thold_posedge$D$CPN$CDN_EQ_1_AN_E_EQ_1 = 1.0,
       tsetup_posedge$E$CPN$CDN_EQ_1 = 1.0,
       thold_posedge$E$CPN$CDN_EQ_1 = 1.0,
       trec$CDN$CPN$D_EQ_1_AN_E_EQ_1 = 1.0,
       trem$CDN$CPN$D_EQ_1_AN_E_EQ_1 = 1.0;

     // path delays
     (negedge CPN *> (QN -: E?D:N_S_XM3_G)) = (tphlh$CPN$QN, tphhl$CPN$QN);
     (negedge CPN *> (Q +: E?D:N_S_XM3_G)) = (tphlh$CPN$Q, tphhl$CPN$Q);
     (negedge CDN *> (QN +: 1'b1)) = (tphlh$CDN$QN, 0);
     (negedge CDN *> (Q -: 1'b1)) = (0, tphhl$CDN$Q);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_E_EQ_1 == 1'b1, negedge D, tsetup_negedge$D$CPN$CDN_EQ_1_AN_E_EQ_1, thold_negedge$D$CPN$CDN_EQ_1_AN_E_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& CDN == 1'b1, negedge E, tsetup_negedge$E$CPN$CDN_EQ_1, thold_negedge$E$CPN$CDN_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_E_EQ_1 == 1'b1, posedge D, tsetup_posedge$D$CPN$CDN_EQ_1_AN_E_EQ_1, thold_posedge$D$CPN$CDN_EQ_1_AN_E_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& CDN == 1'b1, posedge E, tsetup_posedge$E$CPN$CDN_EQ_1, thold_posedge$E$CPN$CDN_EQ_1, NOTIFIER);
     $recrem(posedge CDN, negedge CPN &&& D_EQ_1_AN_E_EQ_1 == 1'b1, trec$CDN$CPN$D_EQ_1_AN_E_EQ_1, trem$CDN$CPN$D_EQ_1_AN_E_EQ_1, NOTIFIER);
     $width(negedge CDN &&& D_EQ_0_AN_E_EQ_0 == 1'b1, tminpwl$CDN$D_EQ_0_AN_E_EQ_0, 0, NOTIFIER);
     $width(posedge CPN &&& CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1 == 1'b1, tminpwh$CPN$CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1, 0, NOTIFIER);
     $width(negedge CPN &&& CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1 == 1'b1, tminpwl$CPN$CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF06ED2 (Q, QN, CDN, CPN, D, E);
input  CDN ;
input  CPN ;
input  D ;
input  E ;
output Q ;
output QN ;
reg NOTIFIER ;

   udp_mux2 (I0_D, N_S_XM3_G, D, E);
   not (I0_CLOCK, CPN);
   not (I0_CLEAR, CDN);
   udp_dff (N_S_XM3_G, I0_D, I0_CLOCK, I0_CLEAR, 1'B0, NOTIFIER);
   not (N_NET0235_XM31_G, N_S_XM3_G);
   not (Q, N_NET0235_XM31_G);
   not (QN, N_S_XM3_G);
   and (CDN_EQ_1_AN_E_EQ_1, CDN, E);
   and (D_EQ_1_AN_E_EQ_1, D, E);
   not (I10_out, D);
   not (I11_out, E);
   and (D_EQ_0_AN_E_EQ_0, I10_out, I11_out);
   not (I13_out, D);
   and (CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1, CDN, I13_out, E);

   specify
     // delay parameters
     specparam
       tphhl$CDN$Q = 1.0,
       tphlh$CDN$QN = 1.0,
       tphlh$CPN$Q = 1.0,
       tphhl$CPN$Q = 1.0,
       tphlh$CPN$QN = 1.0,
       tphhl$CPN$QN = 1.0,
       tminpwl$CDN$D_EQ_0_AN_E_EQ_0 = 1.0,
       tminpwh$CPN$CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1 = 1.0,
       tminpwl$CPN$CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1 = 1.0,
       tsetup_negedge$D$CPN$CDN_EQ_1_AN_E_EQ_1 = 1.0,
       thold_negedge$D$CPN$CDN_EQ_1_AN_E_EQ_1 = 1.0,
       tsetup_negedge$E$CPN$CDN_EQ_1 = 1.0,
       thold_negedge$E$CPN$CDN_EQ_1 = 1.0,
       tsetup_posedge$D$CPN$CDN_EQ_1_AN_E_EQ_1 = 1.0,
       thold_posedge$D$CPN$CDN_EQ_1_AN_E_EQ_1 = 1.0,
       tsetup_posedge$E$CPN$CDN_EQ_1 = 1.0,
       thold_posedge$E$CPN$CDN_EQ_1 = 1.0,
       trec$CDN$CPN$D_EQ_1_AN_E_EQ_1 = 1.0,
       trem$CDN$CPN$D_EQ_1_AN_E_EQ_1 = 1.0;

     // path delays
     (negedge CPN *> (QN -: E?D:N_S_XM3_G)) = (tphlh$CPN$QN, tphhl$CPN$QN);
     (negedge CPN *> (Q +: E?D:N_S_XM3_G)) = (tphlh$CPN$Q, tphhl$CPN$Q);
     (negedge CDN *> (QN +: 1'b1)) = (tphlh$CDN$QN, 0);
     (negedge CDN *> (Q -: 1'b1)) = (0, tphhl$CDN$Q);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_E_EQ_1 == 1'b1, negedge D, tsetup_negedge$D$CPN$CDN_EQ_1_AN_E_EQ_1, thold_negedge$D$CPN$CDN_EQ_1_AN_E_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& CDN == 1'b1, negedge E, tsetup_negedge$E$CPN$CDN_EQ_1, thold_negedge$E$CPN$CDN_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_E_EQ_1 == 1'b1, posedge D, tsetup_posedge$D$CPN$CDN_EQ_1_AN_E_EQ_1, thold_posedge$D$CPN$CDN_EQ_1_AN_E_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& CDN == 1'b1, posedge E, tsetup_posedge$E$CPN$CDN_EQ_1, thold_posedge$E$CPN$CDN_EQ_1, NOTIFIER);
     $recrem(posedge CDN, negedge CPN &&& D_EQ_1_AN_E_EQ_1 == 1'b1, trec$CDN$CPN$D_EQ_1_AN_E_EQ_1, trem$CDN$CPN$D_EQ_1_AN_E_EQ_1, NOTIFIER);
     $width(negedge CDN &&& D_EQ_0_AN_E_EQ_0 == 1'b1, tminpwl$CDN$D_EQ_0_AN_E_EQ_0, 0, NOTIFIER);
     $width(posedge CPN &&& CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1 == 1'b1, tminpwh$CPN$CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1, 0, NOTIFIER);
     $width(negedge CPN &&& CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1 == 1'b1, tminpwl$CPN$CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF06ED4 (Q, QN, CDN, CPN, D, E);
input  CDN ;
input  CPN ;
input  D ;
input  E ;
output Q ;
output QN ;
reg NOTIFIER ;

   udp_mux2 (I0_D, N_S_XM3_G, D, E);
   not (I0_CLOCK, CPN);
   not (I0_CLEAR, CDN);
   udp_dff (N_S_XM3_G, I0_D, I0_CLOCK, I0_CLEAR, 1'B0, NOTIFIER);
   not (N_NET0235_XM31_G, N_S_XM3_G);
   not (Q, N_NET0235_XM31_G);
   not (QN, N_S_XM3_G);
   and (CDN_EQ_1_AN_E_EQ_1, CDN, E);
   and (D_EQ_1_AN_E_EQ_1, D, E);
   not (I10_out, D);
   not (I11_out, E);
   and (D_EQ_0_AN_E_EQ_0, I10_out, I11_out);
   not (I13_out, D);
   and (CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1, CDN, I13_out, E);

   specify
     // delay parameters
     specparam
       tphhl$CDN$Q = 1.0,
       tphlh$CDN$QN = 1.0,
       tphlh$CPN$Q = 1.0,
       tphhl$CPN$Q = 1.0,
       tphlh$CPN$QN = 1.0,
       tphhl$CPN$QN = 1.0,
       tminpwl$CDN$D_EQ_0_AN_E_EQ_0 = 1.0,
       tminpwh$CPN$CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1 = 1.0,
       tminpwl$CPN$CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1 = 1.0,
       tsetup_negedge$D$CPN$CDN_EQ_1_AN_E_EQ_1 = 1.0,
       thold_negedge$D$CPN$CDN_EQ_1_AN_E_EQ_1 = 1.0,
       tsetup_negedge$E$CPN$CDN_EQ_1 = 1.0,
       thold_negedge$E$CPN$CDN_EQ_1 = 1.0,
       tsetup_posedge$D$CPN$CDN_EQ_1_AN_E_EQ_1 = 1.0,
       thold_posedge$D$CPN$CDN_EQ_1_AN_E_EQ_1 = 1.0,
       tsetup_posedge$E$CPN$CDN_EQ_1 = 1.0,
       thold_posedge$E$CPN$CDN_EQ_1 = 1.0,
       trec$CDN$CPN$D_EQ_1_AN_E_EQ_1 = 1.0,
       trem$CDN$CPN$D_EQ_1_AN_E_EQ_1 = 1.0;

     // path delays
     (negedge CPN *> (QN -: E?D:N_S_XM3_G)) = (tphlh$CPN$QN, tphhl$CPN$QN);
     (negedge CPN *> (Q +: E?D:N_S_XM3_G)) = (tphlh$CPN$Q, tphhl$CPN$Q);
     (negedge CDN *> (QN +: 1'b1)) = (tphlh$CDN$QN, 0);
     (negedge CDN *> (Q -: 1'b1)) = (0, tphhl$CDN$Q);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_E_EQ_1 == 1'b1, negedge D, tsetup_negedge$D$CPN$CDN_EQ_1_AN_E_EQ_1, thold_negedge$D$CPN$CDN_EQ_1_AN_E_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& CDN == 1'b1, negedge E, tsetup_negedge$E$CPN$CDN_EQ_1, thold_negedge$E$CPN$CDN_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_E_EQ_1 == 1'b1, posedge D, tsetup_posedge$D$CPN$CDN_EQ_1_AN_E_EQ_1, thold_posedge$D$CPN$CDN_EQ_1_AN_E_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& CDN == 1'b1, posedge E, tsetup_posedge$E$CPN$CDN_EQ_1, thold_posedge$E$CPN$CDN_EQ_1, NOTIFIER);
     $recrem(posedge CDN, negedge CPN &&& D_EQ_1_AN_E_EQ_1 == 1'b1, trec$CDN$CPN$D_EQ_1_AN_E_EQ_1, trem$CDN$CPN$D_EQ_1_AN_E_EQ_1, NOTIFIER);
     $width(negedge CDN &&& D_EQ_0_AN_E_EQ_0 == 1'b1, tminpwl$CDN$D_EQ_0_AN_E_EQ_0, 0, NOTIFIER);
     $width(posedge CPN &&& CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1 == 1'b1, tminpwh$CPN$CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1, 0, NOTIFIER);
     $width(negedge CPN &&& CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1 == 1'b1, tminpwl$CPN$CDN_EQ_1_AN_D_EQ_0_AN_E_EQ_1, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF06HD1 (Q, CDN, CPN, D);
input  CDN ;
input  CPN ;
input  D ;
output Q ;
reg NOTIFIER ;

   not (I0_CLOCK, CPN);
   not (I0_CLEAR, CDN);
   udp_dff (N_S_XM23_G, D, I0_CLOCK, I0_CLEAR, 1'B0, NOTIFIER);
   not (N_NET0130_XM20_D, N_S_XM23_G);
   not (Q, N_NET0130_XM20_D);
   not (I6_out, D);
   and (CDN_EQ_1_AN_D_EQ_0, CDN, I6_out);

   specify
     // delay parameters
     specparam
       tphhl$CDN$Q = 1.0,
       tphlh$CPN$Q = 1.0,
       tphhl$CPN$Q = 1.0,
       tminpwl$CDN$D_EQ_0 = 1.0,
       tminpwh$CPN$CDN_EQ_1_AN_D_EQ_0 = 1.0,
       tminpwl$CPN$CDN_EQ_1_AN_D_EQ_0 = 1.0,
       tsetup_negedge$D$CPN$CDN_EQ_1 = 1.0,
       thold_negedge$D$CPN$CDN_EQ_1 = 1.0,
       tsetup_posedge$D$CPN$CDN_EQ_1 = 1.0,
       thold_posedge$D$CPN$CDN_EQ_1 = 1.0,
       trec$CDN$CPN$D_EQ_1 = 1.0,
       trem$CDN$CPN$D_EQ_1 = 1.0;

     // path delays
     (negedge CPN *> (Q +: D)) = (tphlh$CPN$Q, tphhl$CPN$Q);
     (negedge CDN *> (Q -: 1'b1)) = (0, tphhl$CDN$Q);
     $setuphold(negedge CPN &&& CDN == 1'b1, negedge D, tsetup_negedge$D$CPN$CDN_EQ_1, thold_negedge$D$CPN$CDN_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& CDN == 1'b1, posedge D, tsetup_posedge$D$CPN$CDN_EQ_1, thold_posedge$D$CPN$CDN_EQ_1, NOTIFIER);
     $recrem(posedge CDN, negedge CPN &&& D == 1'b1, trec$CDN$CPN$D_EQ_1, trem$CDN$CPN$D_EQ_1, NOTIFIER);
     $width(negedge CDN &&& D == 1'b0, tminpwl$CDN$D_EQ_0, 0, NOTIFIER);
     $width(posedge CPN &&& CDN_EQ_1_AN_D_EQ_0 == 1'b1, tminpwh$CPN$CDN_EQ_1_AN_D_EQ_0, 0, NOTIFIER);
     $width(negedge CPN &&& CDN_EQ_1_AN_D_EQ_0 == 1'b1, tminpwl$CPN$CDN_EQ_1_AN_D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF06HD2 (Q, CDN, CPN, D);
input  CDN ;
input  CPN ;
input  D ;
output Q ;
reg NOTIFIER ;

   not (I0_CLOCK, CPN);
   not (I0_CLEAR, CDN);
   udp_dff (N_S_XM23_G, D, I0_CLOCK, I0_CLEAR, 1'B0, NOTIFIER);
   not (N_NET0130_XM20_D, N_S_XM23_G);
   not (Q, N_NET0130_XM20_D);
   not (I6_out, D);
   and (CDN_EQ_1_AN_D_EQ_0, CDN, I6_out);

   specify
     // delay parameters
     specparam
       tphhl$CDN$Q = 1.0,
       tphlh$CPN$Q = 1.0,
       tphhl$CPN$Q = 1.0,
       tminpwl$CDN$D_EQ_0 = 1.0,
       tminpwh$CPN$CDN_EQ_1_AN_D_EQ_0 = 1.0,
       tminpwl$CPN$CDN_EQ_1_AN_D_EQ_0 = 1.0,
       tsetup_negedge$D$CPN$CDN_EQ_1 = 1.0,
       thold_negedge$D$CPN$CDN_EQ_1 = 1.0,
       tsetup_posedge$D$CPN$CDN_EQ_1 = 1.0,
       thold_posedge$D$CPN$CDN_EQ_1 = 1.0,
       trec$CDN$CPN$D_EQ_1 = 1.0,
       trem$CDN$CPN$D_EQ_1 = 1.0;

     // path delays
     (negedge CPN *> (Q +: D)) = (tphlh$CPN$Q, tphhl$CPN$Q);
     (negedge CDN *> (Q -: 1'b1)) = (0, tphhl$CDN$Q);
     $setuphold(negedge CPN &&& CDN == 1'b1, negedge D, tsetup_negedge$D$CPN$CDN_EQ_1, thold_negedge$D$CPN$CDN_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& CDN == 1'b1, posedge D, tsetup_posedge$D$CPN$CDN_EQ_1, thold_posedge$D$CPN$CDN_EQ_1, NOTIFIER);
     $recrem(posedge CDN, negedge CPN &&& D == 1'b1, trec$CDN$CPN$D_EQ_1, trem$CDN$CPN$D_EQ_1, NOTIFIER);
     $width(negedge CDN &&& D == 1'b0, tminpwl$CDN$D_EQ_0, 0, NOTIFIER);
     $width(posedge CPN &&& CDN_EQ_1_AN_D_EQ_0 == 1'b1, tminpwh$CPN$CDN_EQ_1_AN_D_EQ_0, 0, NOTIFIER);
     $width(negedge CPN &&& CDN_EQ_1_AN_D_EQ_0 == 1'b1, tminpwl$CPN$CDN_EQ_1_AN_D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF06HD4 (Q, CDN, CPN, D);
input  CDN ;
input  CPN ;
input  D ;
output Q ;
reg NOTIFIER ;

   not (I0_CLOCK, CPN);
   not (I0_CLEAR, CDN);
   udp_dff (N_S_XM23_G, D, I0_CLOCK, I0_CLEAR, 1'B0, NOTIFIER);
   not (N_NET0130_XM20_D, N_S_XM23_G);
   not (Q, N_NET0130_XM20_D);
   not (I6_out, D);
   and (CDN_EQ_1_AN_D_EQ_0, CDN, I6_out);

   specify
     // delay parameters
     specparam
       tphhl$CDN$Q = 1.0,
       tphlh$CPN$Q = 1.0,
       tphhl$CPN$Q = 1.0,
       tminpwl$CDN$D_EQ_0 = 1.0,
       tminpwh$CPN$CDN_EQ_1_AN_D_EQ_0 = 1.0,
       tminpwl$CPN$CDN_EQ_1_AN_D_EQ_0 = 1.0,
       tsetup_negedge$D$CPN$CDN_EQ_1 = 1.0,
       thold_negedge$D$CPN$CDN_EQ_1 = 1.0,
       tsetup_posedge$D$CPN$CDN_EQ_1 = 1.0,
       thold_posedge$D$CPN$CDN_EQ_1 = 1.0,
       trec$CDN$CPN$D_EQ_1 = 1.0,
       trem$CDN$CPN$D_EQ_1 = 1.0;

     // path delays
     (negedge CPN *> (Q +: D)) = (tphlh$CPN$Q, tphhl$CPN$Q);
     (negedge CDN *> (Q -: 1'b1)) = (0, tphhl$CDN$Q);
     $setuphold(negedge CPN &&& CDN == 1'b1, negedge D, tsetup_negedge$D$CPN$CDN_EQ_1, thold_negedge$D$CPN$CDN_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& CDN == 1'b1, posedge D, tsetup_posedge$D$CPN$CDN_EQ_1, thold_posedge$D$CPN$CDN_EQ_1, NOTIFIER);
     $recrem(posedge CDN, negedge CPN &&& D == 1'b1, trec$CDN$CPN$D_EQ_1, trem$CDN$CPN$D_EQ_1, NOTIFIER);
     $width(negedge CDN &&& D == 1'b0, tminpwl$CDN$D_EQ_0, 0, NOTIFIER);
     $width(posedge CPN &&& CDN_EQ_1_AN_D_EQ_0 == 1'b1, tminpwh$CPN$CDN_EQ_1_AN_D_EQ_0, 0, NOTIFIER);
     $width(negedge CPN &&& CDN_EQ_1_AN_D_EQ_0 == 1'b1, tminpwl$CPN$CDN_EQ_1_AN_D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF07D1 (Q, QN, CPN, D, SDN);
input  CPN ;
input  D ;
input  SDN ;
output Q ;
output QN ;
reg NOTIFIER ;

   not (I0_CLOCK, CPN);
   not (I0_SET, SDN);
   udp_dff (N_S_XM21_G, D, I0_CLOCK, 1'B0, I0_SET, NOTIFIER);
   not (N_NET0130_XM18_D, N_S_XM21_G);
   buf (Q, N_S_XM21_G);
   not (QN, N_S_XM21_G);
   not (I8_out, D);
   and (D_EQ_0_AN_SDN_EQ_1, I8_out, SDN);

   specify
     // delay parameters
     specparam
       tphlh$CPN$Q = 1.0,
       tphhl$CPN$Q = 1.0,
       tphlh$CPN$QN = 1.0,
       tphhl$CPN$QN = 1.0,
       tphlh$SDN$Q = 1.0,
       tphhl$SDN$QN = 1.0,
       tminpwh$CPN$D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwl$CPN$D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwl$SDN$D_EQ_0 = 1.0,
       tsetup_negedge$D$CPN$SDN_EQ_1 = 1.0,
       thold_negedge$D$CPN$SDN_EQ_1 = 1.0,
       tsetup_posedge$D$CPN$SDN_EQ_1 = 1.0,
       thold_posedge$D$CPN$SDN_EQ_1 = 1.0,
       trec$SDN$CPN$D_EQ_0 = 1.0,
       trem$SDN$CPN$D_EQ_0 = 1.0;

     // path delays
     (negedge CPN *> (QN -: D)) = (tphlh$CPN$QN, tphhl$CPN$QN);
     (negedge CPN *> (Q +: D)) = (tphlh$CPN$Q, tphhl$CPN$Q);
     (negedge SDN *> (QN -: 1'b1)) = (0, tphhl$SDN$QN);
     (negedge SDN *> (Q +: 1'b1)) = (tphlh$SDN$Q, 0);
     $setuphold(negedge CPN &&& SDN == 1'b1, negedge D, tsetup_negedge$D$CPN$SDN_EQ_1, thold_negedge$D$CPN$SDN_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& SDN == 1'b1, posedge D, tsetup_posedge$D$CPN$SDN_EQ_1, thold_posedge$D$CPN$SDN_EQ_1, NOTIFIER);
     $recrem(posedge SDN, negedge CPN &&& D == 1'b0, trec$SDN$CPN$D_EQ_0, trem$SDN$CPN$D_EQ_0, NOTIFIER);
     $width(posedge CPN &&& D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwh$CPN$D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(negedge CPN &&& D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwl$CPN$D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(negedge SDN &&& D == 1'b0, tminpwl$SDN$D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF07D2 (Q, QN, CPN, D, SDN);
input  CPN ;
input  D ;
input  SDN ;
output Q ;
output QN ;
reg NOTIFIER ;

   not (I0_CLOCK, CPN);
   not (I0_SET, SDN);
   udp_dff (N_S_XM21_G, D, I0_CLOCK, 1'B0, I0_SET, NOTIFIER);
   not (N_NET0130_XM18_D, N_S_XM21_G);
   buf (Q, N_S_XM21_G);
   not (QN, N_S_XM21_G);
   not (I8_out, D);
   and (D_EQ_0_AN_SDN_EQ_1, I8_out, SDN);

   specify
     // delay parameters
     specparam
       tphlh$CPN$Q = 1.0,
       tphhl$CPN$Q = 1.0,
       tphlh$CPN$QN = 1.0,
       tphhl$CPN$QN = 1.0,
       tphlh$SDN$Q = 1.0,
       tphhl$SDN$QN = 1.0,
       tminpwh$CPN$D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwl$CPN$D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwl$SDN$D_EQ_0 = 1.0,
       tsetup_negedge$D$CPN$SDN_EQ_1 = 1.0,
       thold_negedge$D$CPN$SDN_EQ_1 = 1.0,
       tsetup_posedge$D$CPN$SDN_EQ_1 = 1.0,
       thold_posedge$D$CPN$SDN_EQ_1 = 1.0,
       trec$SDN$CPN$D_EQ_0 = 1.0,
       trem$SDN$CPN$D_EQ_0 = 1.0;

     // path delays
     (negedge CPN *> (QN -: D)) = (tphlh$CPN$QN, tphhl$CPN$QN);
     (negedge CPN *> (Q +: D)) = (tphlh$CPN$Q, tphhl$CPN$Q);
     (negedge SDN *> (QN -: 1'b1)) = (0, tphhl$SDN$QN);
     (negedge SDN *> (Q +: 1'b1)) = (tphlh$SDN$Q, 0);
     $setuphold(negedge CPN &&& SDN == 1'b1, negedge D, tsetup_negedge$D$CPN$SDN_EQ_1, thold_negedge$D$CPN$SDN_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& SDN == 1'b1, posedge D, tsetup_posedge$D$CPN$SDN_EQ_1, thold_posedge$D$CPN$SDN_EQ_1, NOTIFIER);
     $recrem(posedge SDN, negedge CPN &&& D == 1'b0, trec$SDN$CPN$D_EQ_0, trem$SDN$CPN$D_EQ_0, NOTIFIER);
     $width(posedge CPN &&& D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwh$CPN$D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(negedge CPN &&& D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwl$CPN$D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(negedge SDN &&& D == 1'b0, tminpwl$SDN$D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF07D4 (Q, QN, CPN, D, SDN);
input  CPN ;
input  D ;
input  SDN ;
output Q ;
output QN ;
reg NOTIFIER ;

   not (I0_CLOCK, CPN);
   not (I0_SET, SDN);
   udp_dff (N_S_XM21_G, D, I0_CLOCK, 1'B0, I0_SET, NOTIFIER);
   not (N_NET0130_XM18_D, N_S_XM21_G);
   buf (Q, N_S_XM21_G);
   not (QN, N_S_XM21_G);
   not (I8_out, D);
   and (D_EQ_0_AN_SDN_EQ_1, I8_out, SDN);

   specify
     // delay parameters
     specparam
       tphlh$CPN$Q = 1.0,
       tphhl$CPN$Q = 1.0,
       tphlh$CPN$QN = 1.0,
       tphhl$CPN$QN = 1.0,
       tphlh$SDN$Q = 1.0,
       tphhl$SDN$QN = 1.0,
       tminpwh$CPN$D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwl$CPN$D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwl$SDN$D_EQ_0 = 1.0,
       tsetup_negedge$D$CPN$SDN_EQ_1 = 1.0,
       thold_negedge$D$CPN$SDN_EQ_1 = 1.0,
       tsetup_posedge$D$CPN$SDN_EQ_1 = 1.0,
       thold_posedge$D$CPN$SDN_EQ_1 = 1.0,
       trec$SDN$CPN$D_EQ_0 = 1.0,
       trem$SDN$CPN$D_EQ_0 = 1.0;

     // path delays
     (negedge CPN *> (QN -: D)) = (tphlh$CPN$QN, tphhl$CPN$QN);
     (negedge CPN *> (Q +: D)) = (tphlh$CPN$Q, tphhl$CPN$Q);
     (negedge SDN *> (QN -: 1'b1)) = (0, tphhl$SDN$QN);
     (negedge SDN *> (Q +: 1'b1)) = (tphlh$SDN$Q, 0);
     $setuphold(negedge CPN &&& SDN == 1'b1, negedge D, tsetup_negedge$D$CPN$SDN_EQ_1, thold_negedge$D$CPN$SDN_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& SDN == 1'b1, posedge D, tsetup_posedge$D$CPN$SDN_EQ_1, thold_posedge$D$CPN$SDN_EQ_1, NOTIFIER);
     $recrem(posedge SDN, negedge CPN &&& D == 1'b0, trec$SDN$CPN$D_EQ_0, trem$SDN$CPN$D_EQ_0, NOTIFIER);
     $width(posedge CPN &&& D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwh$CPN$D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(negedge CPN &&& D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwl$CPN$D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(negedge SDN &&& D == 1'b0, tminpwl$SDN$D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF07HD1 (Q, CPN, D, SDN);
input  CPN ;
input  D ;
input  SDN ;
output Q ;
reg NOTIFIER ;

   not (I0_CLOCK, CPN);
   not (I0_SET, SDN);
   udp_dff (N_S_XM21_G, D, I0_CLOCK, 1'B0, I0_SET, NOTIFIER);
   not (N_NET0130_XM18_D, N_S_XM21_G);
   not (Q, N_NET0130_XM18_D);
   not (I6_out, D);
   and (D_EQ_0_AN_SDN_EQ_1, I6_out, SDN);

   specify
     // delay parameters
     specparam
       tphlh$CPN$Q = 1.0,
       tphhl$CPN$Q = 1.0,
       tphlh$SDN$Q = 1.0,
       tminpwh$CPN$D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwl$CPN$D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwl$SDN$D_EQ_0 = 1.0,
       tsetup_negedge$D$CPN$SDN_EQ_1 = 1.0,
       thold_negedge$D$CPN$SDN_EQ_1 = 1.0,
       tsetup_posedge$D$CPN$SDN_EQ_1 = 1.0,
       thold_posedge$D$CPN$SDN_EQ_1 = 1.0,
       trec$SDN$CPN$D_EQ_0 = 1.0,
       trem$SDN$CPN$D_EQ_0 = 1.0;

     // path delays
     (negedge CPN *> (Q +: D)) = (tphlh$CPN$Q, tphhl$CPN$Q);
     (negedge SDN *> (Q +: 1'b1)) = (tphlh$SDN$Q, 0);
     $setuphold(negedge CPN &&& SDN == 1'b1, negedge D, tsetup_negedge$D$CPN$SDN_EQ_1, thold_negedge$D$CPN$SDN_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& SDN == 1'b1, posedge D, tsetup_posedge$D$CPN$SDN_EQ_1, thold_posedge$D$CPN$SDN_EQ_1, NOTIFIER);
     $recrem(posedge SDN, negedge CPN &&& D == 1'b0, trec$SDN$CPN$D_EQ_0, trem$SDN$CPN$D_EQ_0, NOTIFIER);
     $width(posedge CPN &&& D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwh$CPN$D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(negedge CPN &&& D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwl$CPN$D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(negedge SDN &&& D == 1'b0, tminpwl$SDN$D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF07HD2 (Q, CPN, D, SDN);
input  CPN ;
input  D ;
input  SDN ;
output Q ;
reg NOTIFIER ;

   not (I0_CLOCK, CPN);
   not (I0_SET, SDN);
   udp_dff (N_S_XM21_G, D, I0_CLOCK, 1'B0, I0_SET, NOTIFIER);
   not (N_NET0130_XM18_D, N_S_XM21_G);
   not (Q, N_NET0130_XM18_D);
   not (I6_out, D);
   and (D_EQ_0_AN_SDN_EQ_1, I6_out, SDN);

   specify
     // delay parameters
     specparam
       tphlh$CPN$Q = 1.0,
       tphhl$CPN$Q = 1.0,
       tphlh$SDN$Q = 1.0,
       tminpwh$CPN$D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwl$CPN$D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwl$SDN$D_EQ_0 = 1.0,
       tsetup_negedge$D$CPN$SDN_EQ_1 = 1.0,
       thold_negedge$D$CPN$SDN_EQ_1 = 1.0,
       tsetup_posedge$D$CPN$SDN_EQ_1 = 1.0,
       thold_posedge$D$CPN$SDN_EQ_1 = 1.0,
       trec$SDN$CPN$D_EQ_0 = 1.0,
       trem$SDN$CPN$D_EQ_0 = 1.0;

     // path delays
     (negedge CPN *> (Q +: D)) = (tphlh$CPN$Q, tphhl$CPN$Q);
     (negedge SDN *> (Q +: 1'b1)) = (tphlh$SDN$Q, 0);
     $setuphold(negedge CPN &&& SDN == 1'b1, negedge D, tsetup_negedge$D$CPN$SDN_EQ_1, thold_negedge$D$CPN$SDN_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& SDN == 1'b1, posedge D, tsetup_posedge$D$CPN$SDN_EQ_1, thold_posedge$D$CPN$SDN_EQ_1, NOTIFIER);
     $recrem(posedge SDN, negedge CPN &&& D == 1'b0, trec$SDN$CPN$D_EQ_0, trem$SDN$CPN$D_EQ_0, NOTIFIER);
     $width(posedge CPN &&& D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwh$CPN$D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(negedge CPN &&& D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwl$CPN$D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(negedge SDN &&& D == 1'b0, tminpwl$SDN$D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF07HD4 (Q, CPN, D, SDN);
input  CPN ;
input  D ;
input  SDN ;
output Q ;
reg NOTIFIER ;

   not (I0_CLOCK, CPN);
   not (I0_SET, SDN);
   udp_dff (N_S_XM21_G, D, I0_CLOCK, 1'B0, I0_SET, NOTIFIER);
   not (N_NET0130_XM18_D, N_S_XM21_G);
   not (Q, N_NET0130_XM18_D);
   not (I6_out, D);
   and (D_EQ_0_AN_SDN_EQ_1, I6_out, SDN);

   specify
     // delay parameters
     specparam
       tphlh$CPN$Q = 1.0,
       tphhl$CPN$Q = 1.0,
       tphlh$SDN$Q = 1.0,
       tminpwh$CPN$D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwl$CPN$D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwl$SDN$D_EQ_0 = 1.0,
       tsetup_negedge$D$CPN$SDN_EQ_1 = 1.0,
       thold_negedge$D$CPN$SDN_EQ_1 = 1.0,
       tsetup_posedge$D$CPN$SDN_EQ_1 = 1.0,
       thold_posedge$D$CPN$SDN_EQ_1 = 1.0,
       trec$SDN$CPN$D_EQ_0 = 1.0,
       trem$SDN$CPN$D_EQ_0 = 1.0;

     // path delays
     (negedge CPN *> (Q +: D)) = (tphlh$CPN$Q, tphhl$CPN$Q);
     (negedge SDN *> (Q +: 1'b1)) = (tphlh$SDN$Q, 0);
     $setuphold(negedge CPN &&& SDN == 1'b1, negedge D, tsetup_negedge$D$CPN$SDN_EQ_1, thold_negedge$D$CPN$SDN_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& SDN == 1'b1, posedge D, tsetup_posedge$D$CPN$SDN_EQ_1, thold_posedge$D$CPN$SDN_EQ_1, NOTIFIER);
     $recrem(posedge SDN, negedge CPN &&& D == 1'b0, trec$SDN$CPN$D_EQ_0, trem$SDN$CPN$D_EQ_0, NOTIFIER);
     $width(posedge CPN &&& D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwh$CPN$D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(negedge CPN &&& D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwl$CPN$D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(negedge SDN &&& D == 1'b0, tminpwl$SDN$D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF08D1 (Q, QN, CDN, CPN, D, SDN);
input  CDN ;
input  CPN ;
input  D ;
input  SDN ;
output Q ;
output QN ;
reg NOTIFIER ;

   not (I0_CLOCK, CPN);
   not (I0_CLEAR, CDN);
   not (I0_SET, SDN);
   udp_dff (N_S_XM25_G, D, I0_CLOCK, I0_CLEAR, I0_SET, NOTIFIER);
   not (N_NET0130_XM22_D, N_S_XM25_G);
   not (Q, N_NET0130_XM22_D);
   buf (QN, N_NET0130_XM22_D);
   not (I9_out, D);
   and (CDN_EQ_1_AN_D_EQ_0, CDN, I9_out);
   and (CDN_EQ_1_AN_SDN_EQ_1, CDN, SDN);
   and (D_EQ_1_AN_SDN_EQ_1, D, SDN);
   not (I13_out, D);
   and (D_EQ_0_AN_SDN_EQ_1, I13_out, SDN);
   not (I15_out, D);
   and (CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1, CDN, I15_out, SDN);
   not (I18_out, CDN);
   not (I19_out, D);
   and (CDN_EQ_0_AN_D_EQ_0, I18_out, I19_out);

   specify
     // delay parameters
     specparam
       tphhl$CDN$Q = 1.0,
       tphlh$CDN$QN = 1.0,
       tphlh$CPN$Q = 1.0,
       tphhl$CPN$Q = 1.0,
       tphlh$CPN$QN = 1.0,
       tphhl$CPN$QN = 1.0,
       tplhl$SDN$Q = 1.0,
       tphlh$SDN$Q = 1.0,
       tpllh$SDN$QN = 1.0,
       tphhl$SDN$QN = 1.0,
       tminpwl$CDN$D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwh$CPN$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwl$CPN$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwl$SDN$CDN_EQ_0_AN_D_EQ_0 = 1.0,
       tsetup_negedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       thold_negedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       tsetup_posedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       thold_posedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       trec$CDN$CPN$D_EQ_1_AN_SDN_EQ_1 = 1.0,
       trem$CDN$CPN$D_EQ_1_AN_SDN_EQ_1 = 1.0,
       trec$CDN$SDN$D_EQ_0 = 1.0,
       trec$SDN$CPN$CDN_EQ_1_AN_D_EQ_0 = 1.0,
       trem$SDN$CPN$CDN_EQ_1_AN_D_EQ_0 = 1.0;

     // path delays
     (negedge CPN *> (QN -: D)) = (tphlh$CPN$QN, tphhl$CPN$QN);
     (negedge CPN *> (Q +: D)) = (tphlh$CPN$Q, tphhl$CPN$Q);
     (negedge SDN *> (QN -: 1'b1)) = (tpllh$SDN$QN, tphhl$SDN$QN);
     (negedge SDN *> (Q +: 1'b1)) = (tphlh$SDN$Q, tplhl$SDN$Q);
     (negedge CDN *> (QN +: 1'b1)) = (tphlh$CDN$QN, 0);
     (negedge CDN *> (Q -: 1'b1)) = (0, tphhl$CDN$Q);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_SDN_EQ_1 == 1'b1, negedge D, tsetup_negedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1, thold_negedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_SDN_EQ_1 == 1'b1, posedge D, tsetup_posedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1, thold_posedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1, NOTIFIER);
     $recrem(posedge CDN, negedge CPN &&& D_EQ_1_AN_SDN_EQ_1 == 1'b1, trec$CDN$CPN$D_EQ_1_AN_SDN_EQ_1, trem$CDN$CPN$D_EQ_1_AN_SDN_EQ_1, NOTIFIER);
     $recovery(posedge CDN, posedge SDN &&& D == 1'b0, trec$CDN$SDN$D_EQ_0, NOTIFIER);
     $recrem(posedge SDN, negedge CPN &&& CDN_EQ_1_AN_D_EQ_0 == 1'b1, trec$SDN$CPN$CDN_EQ_1_AN_D_EQ_0, trem$SDN$CPN$CDN_EQ_1_AN_D_EQ_0, NOTIFIER);
     $width(negedge CDN &&& D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwl$CDN$D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(posedge CPN &&& CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwh$CPN$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(negedge CPN &&& CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwl$CPN$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(negedge SDN &&& CDN_EQ_0_AN_D_EQ_0 == 1'b1, tminpwl$SDN$CDN_EQ_0_AN_D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF08D2 (Q, QN, CDN, CPN, D, SDN);
input  CDN ;
input  CPN ;
input  D ;
input  SDN ;
output Q ;
output QN ;
reg NOTIFIER ;

   not (I0_CLOCK, CPN);
   not (I0_CLEAR, CDN);
   not (I0_SET, SDN);
   udp_dff (N_S_XM25_G, D, I0_CLOCK, I0_CLEAR, I0_SET, NOTIFIER);
   not (N_NET0130_XM22_D, N_S_XM25_G);
   not (Q, N_NET0130_XM22_D);
   buf (QN, N_NET0130_XM22_D);
   not (I9_out, D);
   and (CDN_EQ_1_AN_D_EQ_0, CDN, I9_out);
   and (CDN_EQ_1_AN_SDN_EQ_1, CDN, SDN);
   and (D_EQ_1_AN_SDN_EQ_1, D, SDN);
   not (I13_out, D);
   and (D_EQ_0_AN_SDN_EQ_1, I13_out, SDN);
   not (I15_out, D);
   and (CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1, CDN, I15_out, SDN);
   not (I18_out, CDN);
   not (I19_out, D);
   and (CDN_EQ_0_AN_D_EQ_0, I18_out, I19_out);

   specify
     // delay parameters
     specparam
       tphhl$CDN$Q = 1.0,
       tphlh$CDN$QN = 1.0,
       tphlh$CPN$Q = 1.0,
       tphhl$CPN$Q = 1.0,
       tphlh$CPN$QN = 1.0,
       tphhl$CPN$QN = 1.0,
       tplhl$SDN$Q = 1.0,
       tphlh$SDN$Q = 1.0,
       tpllh$SDN$QN = 1.0,
       tphhl$SDN$QN = 1.0,
       tminpwl$CDN$D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwh$CPN$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwl$CPN$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwl$SDN$CDN_EQ_0_AN_D_EQ_0 = 1.0,
       tsetup_negedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       thold_negedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       tsetup_posedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       thold_posedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       trec$CDN$CPN$D_EQ_1_AN_SDN_EQ_1 = 1.0,
       trem$CDN$CPN$D_EQ_1_AN_SDN_EQ_1 = 1.0,
       trec$CDN$SDN$D_EQ_0 = 1.0,
       trec$SDN$CPN$CDN_EQ_1_AN_D_EQ_0 = 1.0,
       trem$SDN$CPN$CDN_EQ_1_AN_D_EQ_0 = 1.0;

     // path delays
     (negedge CPN *> (QN -: D)) = (tphlh$CPN$QN, tphhl$CPN$QN);
     (negedge CPN *> (Q +: D)) = (tphlh$CPN$Q, tphhl$CPN$Q);
     (negedge SDN *> (QN -: 1'b1)) = (tpllh$SDN$QN, tphhl$SDN$QN);
     (negedge SDN *> (Q +: 1'b1)) = (tphlh$SDN$Q, tplhl$SDN$Q);
     (negedge CDN *> (QN +: 1'b1)) = (tphlh$CDN$QN, 0);
     (negedge CDN *> (Q -: 1'b1)) = (0, tphhl$CDN$Q);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_SDN_EQ_1 == 1'b1, negedge D, tsetup_negedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1, thold_negedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_SDN_EQ_1 == 1'b1, posedge D, tsetup_posedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1, thold_posedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1, NOTIFIER);
     $recrem(posedge CDN, negedge CPN &&& D_EQ_1_AN_SDN_EQ_1 == 1'b1, trec$CDN$CPN$D_EQ_1_AN_SDN_EQ_1, trem$CDN$CPN$D_EQ_1_AN_SDN_EQ_1, NOTIFIER);
     $recovery(posedge CDN, posedge SDN &&& D == 1'b0, trec$CDN$SDN$D_EQ_0, NOTIFIER);
     $recrem(posedge SDN, negedge CPN &&& CDN_EQ_1_AN_D_EQ_0 == 1'b1, trec$SDN$CPN$CDN_EQ_1_AN_D_EQ_0, trem$SDN$CPN$CDN_EQ_1_AN_D_EQ_0, NOTIFIER);
     $width(negedge CDN &&& D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwl$CDN$D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(posedge CPN &&& CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwh$CPN$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(negedge CPN &&& CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwl$CPN$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(negedge SDN &&& CDN_EQ_0_AN_D_EQ_0 == 1'b1, tminpwl$SDN$CDN_EQ_0_AN_D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DF08D4 (Q, QN, CDN, CPN, D, SDN);
input  CDN ;
input  CPN ;
input  D ;
input  SDN ;
output Q ;
output QN ;
reg NOTIFIER ;

   not (I0_CLOCK, CPN);
   not (I0_CLEAR, CDN);
   not (I0_SET, SDN);
   udp_dff (N_S_XM25_G, D, I0_CLOCK, I0_CLEAR, I0_SET, NOTIFIER);
   not (N_NET0130_XM22_D, N_S_XM25_G);
   not (Q, N_NET0130_XM22_D);
   buf (QN, N_NET0130_XM22_D);
   not (I9_out, D);
   and (CDN_EQ_1_AN_D_EQ_0, CDN, I9_out);
   and (CDN_EQ_1_AN_SDN_EQ_1, CDN, SDN);
   and (D_EQ_1_AN_SDN_EQ_1, D, SDN);
   not (I13_out, D);
   and (D_EQ_0_AN_SDN_EQ_1, I13_out, SDN);
   not (I15_out, D);
   and (CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1, CDN, I15_out, SDN);
   not (I18_out, CDN);
   not (I19_out, D);
   and (CDN_EQ_0_AN_D_EQ_0, I18_out, I19_out);

   specify
     // delay parameters
     specparam
       tphhl$CDN$Q = 1.0,
       tphlh$CDN$QN = 1.0,
       tphlh$CPN$Q = 1.0,
       tphhl$CPN$Q = 1.0,
       tphlh$CPN$QN = 1.0,
       tphhl$CPN$QN = 1.0,
       tplhl$SDN$Q = 1.0,
       tphlh$SDN$Q = 1.0,
       tpllh$SDN$QN = 1.0,
       tphhl$SDN$QN = 1.0,
       tminpwl$CDN$D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwh$CPN$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwl$CPN$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwl$SDN$CDN_EQ_0_AN_D_EQ_0 = 1.0,
       tsetup_negedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       thold_negedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       tsetup_posedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       thold_posedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       trec$CDN$CPN$D_EQ_1_AN_SDN_EQ_1 = 1.0,
       trem$CDN$CPN$D_EQ_1_AN_SDN_EQ_1 = 1.0,
       trec$CDN$SDN$D_EQ_0 = 1.0,
       trec$SDN$CPN$CDN_EQ_1_AN_D_EQ_0 = 1.0,
       trem$SDN$CPN$CDN_EQ_1_AN_D_EQ_0 = 1.0;

     // path delays
     (negedge CPN *> (QN -: D)) = (tphlh$CPN$QN, tphhl$CPN$QN);
     (negedge CPN *> (Q +: D)) = (tphlh$CPN$Q, tphhl$CPN$Q);
     (negedge SDN *> (QN -: 1'b1)) = (tpllh$SDN$QN, tphhl$SDN$QN);
     (negedge SDN *> (Q +: 1'b1)) = (tphlh$SDN$Q, tplhl$SDN$Q);
     (negedge CDN *> (QN +: 1'b1)) = (tphlh$CDN$QN, 0);
     (negedge CDN *> (Q -: 1'b1)) = (0, tphhl$CDN$Q);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_SDN_EQ_1 == 1'b1, negedge D, tsetup_negedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1, thold_negedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_SDN_EQ_1 == 1'b1, posedge D, tsetup_posedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1, thold_posedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1, NOTIFIER);
     $recrem(posedge CDN, negedge CPN &&& D_EQ_1_AN_SDN_EQ_1 == 1'b1, trec$CDN$CPN$D_EQ_1_AN_SDN_EQ_1, trem$CDN$CPN$D_EQ_1_AN_SDN_EQ_1, NOTIFIER);
     $recovery(posedge CDN, posedge SDN &&& D == 1'b0, trec$CDN$SDN$D_EQ_0, NOTIFIER);
     $recrem(posedge SDN, negedge CPN &&& CDN_EQ_1_AN_D_EQ_0 == 1'b1, trec$SDN$CPN$CDN_EQ_1_AN_D_EQ_0, trem$SDN$CPN$CDN_EQ_1_AN_D_EQ_0, NOTIFIER);
     $width(negedge CDN &&& D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwl$CDN$D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(posedge CPN &&& CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwh$CPN$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(negedge CPN &&& CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwl$CPN$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(negedge SDN &&& CDN_EQ_0_AN_D_EQ_0 == 1'b1, tminpwl$SDN$CDN_EQ_0_AN_D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DL01D1 (Z, I);
input  I ;
output Z ;

   buf (Z, I);

   specify
     // delay parameters
     specparam
       tpllh$I$Z = 1.0,
       tphhl$I$Z = 1.0;

     // path delays
     (I *> Z) = (tpllh$I$Z, tphhl$I$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DL02D1 (Z, I);
input  I ;
output Z ;

   buf (Z, I);

   specify
     // delay parameters
     specparam
       tpllh$I$Z = 1.0,
       tphhl$I$Z = 1.0;

     // path delays
     (I *> Z) = (tpllh$I$Z, tphhl$I$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DL03D1 (Z, I);
input  I ;
output Z ;

   buf (Z, I);

   specify
     // delay parameters
     specparam
       tpllh$I$Z = 1.0,
       tphhl$I$Z = 1.0;

     // path delays
     (I *> Z) = (tpllh$I$Z, tphhl$I$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DL04D1 (Z, I);
input  I ;
output Z ;

   buf (Z, I);

   specify
     // delay parameters
     specparam
       tpllh$I$Z = 1.0,
       tphhl$I$Z = 1.0;

     // path delays
     (I *> Z) = (tpllh$I$Z, tphhl$I$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DT01D1 (Q, QN, D, E);
input  D ;
input  E ;
output Q ;
output QN ;
reg NOTIFIER ;

   udp_tlat (N_M_XM9_G, D, E, 1'B0, 1'B0, NOTIFIER);
   not (N_NET0208_XM6_D, N_M_XM9_G);
   buf (Q, N_M_XM9_G);
   not (QN, N_M_XM9_G);

   specify
     // delay parameters
     specparam
       tpllh$D$Q = 1.0,
       tphhl$D$Q = 1.0,
       tplhl$D$QN = 1.0,
       tphlh$D$QN = 1.0,
       tpllh$E$Q = 1.0,
       tplhl$E$Q = 1.0,
       tpllh$E$QN = 1.0,
       tplhl$E$QN = 1.0,
       tminpwh$E$D_EQ_0 = 1.0,
       tsetup_negedge$D$E = 1.0,
       thold_negedge$D$E = 1.0,
       tsetup_posedge$D$E = 1.0,
       thold_posedge$D$E = 1.0;

     // path delays
     (posedge E *> (QN -: D)) = (tpllh$E$QN, tplhl$E$QN);
     (posedge E *> (Q +: D)) = (tpllh$E$Q, tplhl$E$Q);
     (D *> QN) = (tphlh$D$QN, tplhl$D$QN);
     (D *> Q) = (tpllh$D$Q, tphhl$D$Q);
     $setuphold(negedge E, negedge D, tsetup_negedge$D$E, thold_negedge$D$E, NOTIFIER);
     $setuphold(negedge E, posedge D, tsetup_posedge$D$E, thold_posedge$D$E, NOTIFIER);
     $width(posedge E &&& D == 1'b0, tminpwh$E$D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DT02D1 (Q, QN, CDN, D, E);
input  CDN ;
input  D ;
input  E ;
output Q ;
output QN ;
reg NOTIFIER ;

   not (I0_CLEAR, CDN);
   udp_tlat (N_M_XM11_G, D, E, I0_CLEAR, 1'B0, NOTIFIER);
   not (N_NET53_XM5_D, N_M_XM11_G);
   buf (Q, N_M_XM11_G);
   not (QN, N_M_XM11_G);
   not (I7_out, D);
   and (CDN_EQ_1_AN_D_EQ_0, CDN, I7_out);

   specify
     // delay parameters
     specparam
       tpllh$D$Q = 1.0,
       tphhl$D$Q = 1.0,
       tplhl$D$QN = 1.0,
       tphlh$D$QN = 1.0,
       tpllh$CDN$Q = 1.0,
       tphhl$CDN$Q = 1.0,
       tplhl$CDN$QN = 1.0,
       tphlh$CDN$QN = 1.0,
       tpllh$E$Q = 1.0,
       tplhl$E$Q = 1.0,
       tpllh$E$QN = 1.0,
       tplhl$E$QN = 1.0,
       tminpwl$CDN$D_EQ_0 = 1.0,
       tminpwh$E$CDN_EQ_1_AN_D_EQ_0 = 1.0,
       tsetup_negedge$D$E$CDN_EQ_1 = 1.0,
       thold_negedge$D$E$CDN_EQ_1 = 1.0,
       tsetup_posedge$D$E$CDN_EQ_1 = 1.0,
       thold_posedge$D$E$CDN_EQ_1 = 1.0,
       trec$CDN$E$D_EQ_1 = 1.0,
       trem$CDN$E$D_EQ_1 = 1.0;

     // path delays
     (posedge E *> (QN -: D)) = (tpllh$E$QN, tplhl$E$QN);
     (posedge E *> (Q +: D)) = (tpllh$E$Q, tplhl$E$Q);
     (D *> QN) = (tphlh$D$QN, tplhl$D$QN);
     (D *> Q) = (tpllh$D$Q, tphhl$D$Q);
     (negedge CDN *> (QN -: 1'b0)) = (tphlh$CDN$QN, tplhl$CDN$QN);
     (negedge CDN *> (Q +: 1'b0)) = (tpllh$CDN$Q, tphhl$CDN$Q);
     $setuphold(negedge E &&& CDN == 1'b1, negedge D, tsetup_negedge$D$E$CDN_EQ_1, thold_negedge$D$E$CDN_EQ_1, NOTIFIER);
     $setuphold(negedge E &&& CDN == 1'b1, posedge D, tsetup_posedge$D$E$CDN_EQ_1, thold_posedge$D$E$CDN_EQ_1, NOTIFIER);
     $recrem(posedge CDN, negedge E &&& D == 1'b1, trec$CDN$E$D_EQ_1, trem$CDN$E$D_EQ_1, NOTIFIER);
     $width(negedge CDN &&& D == 1'b0, tminpwl$CDN$D_EQ_0, 0, NOTIFIER);
     $width(posedge E &&& CDN_EQ_1_AN_D_EQ_0 == 1'b1, tminpwh$E$CDN_EQ_1_AN_D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_DT03D1 (Q, QN, D, E, SDN);
input  D ;
input  E ;
input  SDN ;
output Q ;
output QN ;
reg NOTIFIER ;

   not (I0_SET, SDN);
   udp_tlat (N_M_XM13_G, D, E, 1'B0, I0_SET, NOTIFIER);
   not (N_NET0208_XM10_D, N_M_XM13_G);
   buf (Q, N_M_XM13_G);
   not (QN, N_M_XM13_G);
   not (I7_out, D);
   and (D_EQ_0_AN_SDN_EQ_1, I7_out, SDN);

   specify
     // delay parameters
     specparam
       tpllh$D$Q = 1.0,
       tphhl$D$Q = 1.0,
       tplhl$D$QN = 1.0,
       tphlh$D$QN = 1.0,
       tpllh$E$Q = 1.0,
       tplhl$E$Q = 1.0,
       tpllh$E$QN = 1.0,
       tplhl$E$QN = 1.0,
       tplhl$SDN$Q = 1.0,
       tphlh$SDN$Q = 1.0,
       tpllh$SDN$QN = 1.0,
       tphhl$SDN$QN = 1.0,
       tminpwh$E$D_EQ_0_AN_SDN_EQ_1 = 1.0,
       tminpwl$SDN$D_EQ_0 = 1.0,
       tsetup_negedge$D$E$SDN_EQ_1 = 1.0,
       thold_negedge$D$E$SDN_EQ_1 = 1.0,
       tsetup_posedge$D$E$SDN_EQ_1 = 1.0,
       thold_posedge$D$E$SDN_EQ_1 = 1.0,
       trec$SDN$E$D_EQ_0 = 1.0,
       trem$SDN$E$D_EQ_0 = 1.0;

     // path delays
     (posedge E *> (QN -: D)) = (tpllh$E$QN, tplhl$E$QN);
     (posedge E *> (Q +: D)) = (tpllh$E$Q, tplhl$E$Q);
     (negedge SDN *> (QN -: 1'b1)) = (tpllh$SDN$QN, tphhl$SDN$QN);
     (negedge SDN *> (Q +: 1'b1)) = (tphlh$SDN$Q, tplhl$SDN$Q);
     (D *> QN) = (tphlh$D$QN, tplhl$D$QN);
     (D *> Q) = (tpllh$D$Q, tphhl$D$Q);
     $setuphold(negedge E &&& SDN == 1'b1, negedge D, tsetup_negedge$D$E$SDN_EQ_1, thold_negedge$D$E$SDN_EQ_1, NOTIFIER);
     $setuphold(negedge E &&& SDN == 1'b1, posedge D, tsetup_posedge$D$E$SDN_EQ_1, thold_posedge$D$E$SDN_EQ_1, NOTIFIER);
     $recrem(posedge SDN, negedge E &&& D == 1'b0, trec$SDN$E$D_EQ_0, trem$SDN$E$D_EQ_0, NOTIFIER);
     $width(posedge E &&& D_EQ_0_AN_SDN_EQ_1 == 1'b1, tminpwh$E$D_EQ_0_AN_SDN_EQ_1, 0, NOTIFIER);
     $width(negedge SDN &&& D == 1'b0, tminpwl$SDN$D_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_FA01D1 (CO, S, A, B, CI);
input  A ;
input  B ;
input  CI ;
output CO ;
output S ;

   and (I0_out, A, B);
   and (I1_out, B, CI);
   and (I3_out, CI, A);
   or  (CO, I0_out, I1_out, I3_out);
   xor (I5_out, A, B);
   xor (S, I5_out, CI);

   specify
     // delay parameters
   /*  specparam
       tpllh$A$S = 1.0,
       tplhl$A$S = 1.0,
       tphlh$A$S = 1.0,
       tphhl$A$S = 1.0,
       tpllh$A$CO = 1.0,
       tphhl$A$CO = 1.0,
       tpllh$B$S = 1.0,
       tplhl$B$S = 1.0,
       tphlh$B$S = 1.0,
       tphhl$B$S = 1.0,
       tpllh$B$CO = 1.0,
       tphhl$B$CO = 1.0,
       tpllh$CI$S = 1.0,
       tplhl$CI$S = 1.0,
       tphlh$CI$S = 1.0,
       tphhl$CI$S = 1.0,
       tpllh$CI$CO = 1.0,
       tphhl$CI$CO = 1.0,
       tpllh$A$S$B_EQ_1_AN_CI_EQ_1 = 1.0,
       tphhl$A$S$B_EQ_1_AN_CI_EQ_1 = 1.0,
       tpllh$A$S$B_EQ_0_AN_CI_EQ_0 = 1.0,
       tphhl$A$S$B_EQ_0_AN_CI_EQ_0 = 1.0,
       tplhl$A$S$B_EQ_1_AN_CI_EQ_0 = 1.0,
       tphlh$A$S$B_EQ_1_AN_CI_EQ_0 = 1.0,
       tplhl$A$S$B_EQ_0_AN_CI_EQ_1 = 1.0,
       tphlh$A$S$B_EQ_0_AN_CI_EQ_1 = 1.0,
       tpllh$A$CO$B_EQ_1_AN_CI_EQ_0 = 1.0,
       tphhl$A$CO$B_EQ_1_AN_CI_EQ_0 = 1.0,
       tpllh$A$CO$B_EQ_0_AN_CI_EQ_1 = 1.0,
       tphhl$A$CO$B_EQ_0_AN_CI_EQ_1 = 1.0,
       tpllh$B$S$A_EQ_1_AN_CI_EQ_1 = 1.0,
       tphhl$B$S$A_EQ_1_AN_CI_EQ_1 = 1.0,
       tpllh$B$S$A_EQ_0_AN_CI_EQ_0 = 1.0,
       tphhl$B$S$A_EQ_0_AN_CI_EQ_0 = 1.0,
       tplhl$B$S$A_EQ_0_AN_CI_EQ_1 = 1.0,
       tphlh$B$S$A_EQ_0_AN_CI_EQ_1 = 1.0,
       tplhl$B$S$A_EQ_1_AN_CI_EQ_0 = 1.0,
       tphlh$B$S$A_EQ_1_AN_CI_EQ_0 = 1.0,
       tpllh$B$CO$A_EQ_1_AN_CI_EQ_0 = 1.0,
       tphhl$B$CO$A_EQ_1_AN_CI_EQ_0 = 1.0,
       tpllh$B$CO$A_EQ_0_AN_CI_EQ_1 = 1.0,
       tphhl$B$CO$A_EQ_0_AN_CI_EQ_1 = 1.0,
       tpllh$CI$S$A_EQ_1_AN_B_EQ_1 = 1.0,
       tphhl$CI$S$A_EQ_1_AN_B_EQ_1 = 1.0,
       tpllh$CI$S$A_EQ_0_AN_B_EQ_0 = 1.0,
       tphhl$CI$S$A_EQ_0_AN_B_EQ_0 = 1.0,
       tplhl$CI$S$A_EQ_1_AN_B_EQ_0 = 1.0,
       tphlh$CI$S$A_EQ_1_AN_B_EQ_0 = 1.0,
       tplhl$CI$S$A_EQ_0_AN_B_EQ_1 = 1.0,
       tphlh$CI$S$A_EQ_0_AN_B_EQ_1 = 1.0,
       tpllh$CI$CO$A_EQ_1_AN_B_EQ_0 = 1.0,
       tphhl$CI$CO$A_EQ_1_AN_B_EQ_0 = 1.0,
       tpllh$CI$CO$A_EQ_0_AN_B_EQ_1 = 1.0,
       tphhl$CI$CO$A_EQ_0_AN_B_EQ_1 = 1.0;

     // path delays
     if (A == 1'b1 && B == 1'b1)
       (CI *> S) = (tpllh$CI$S$A_EQ_1_AN_B_EQ_1, tphhl$CI$S$A_EQ_1_AN_B_EQ_1);
     if (A == 1'b1 && B == 1'b0)
       (CI *> S) = (tphlh$CI$S$A_EQ_1_AN_B_EQ_0, tplhl$CI$S$A_EQ_1_AN_B_EQ_0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> S) = (tphlh$CI$S$A_EQ_0_AN_B_EQ_1, tplhl$CI$S$A_EQ_0_AN_B_EQ_1);
     if (A == 1'b0 && B == 1'b0)
       (CI *> S) = (tpllh$CI$S$A_EQ_0_AN_B_EQ_0, tphhl$CI$S$A_EQ_0_AN_B_EQ_0);
     ifnone
       (CI *> S) = (tpllh$CI$S,tplhl$CI$S);

     if (A == 1'b1 && B == 1'b0)
       (CI *> CO) = (tpllh$CI$CO$A_EQ_1_AN_B_EQ_0, tphhl$CI$CO$A_EQ_1_AN_B_EQ_0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> CO) = (tpllh$CI$CO$A_EQ_0_AN_B_EQ_1, tphhl$CI$CO$A_EQ_0_AN_B_EQ_1);
     ifnone
       (CI *> CO) = (tpllh$CI$CO,tphhl$CI$CO);

     if (A == 1'b1 && CI == 1'b1)
       (B *> S) = (tpllh$B$S$A_EQ_1_AN_CI_EQ_1, tphhl$B$S$A_EQ_1_AN_CI_EQ_1);
     if (A == 1'b1 && CI == 1'b0)
       (B *> S) = (tphlh$B$S$A_EQ_1_AN_CI_EQ_0, tplhl$B$S$A_EQ_1_AN_CI_EQ_0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> S) = (tphlh$B$S$A_EQ_0_AN_CI_EQ_1, tplhl$B$S$A_EQ_0_AN_CI_EQ_1);
     if (A == 1'b0 && CI == 1'b0)
       (B *> S) = (tpllh$B$S$A_EQ_0_AN_CI_EQ_0, tphhl$B$S$A_EQ_0_AN_CI_EQ_0);
     ifnone
       (B *> S) = (tpllh$B$S,tplhl$B$S);

     if (A == 1'b1 && CI == 1'b0)
       (B *> CO) = (tpllh$B$CO$A_EQ_1_AN_CI_EQ_0, tphhl$B$CO$A_EQ_1_AN_CI_EQ_0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> CO) = (tpllh$B$CO$A_EQ_0_AN_CI_EQ_1, tphhl$B$CO$A_EQ_0_AN_CI_EQ_1);
     ifnone
       (B *> CO) = (tpllh$B$CO,tphhl$B$CO);

     if (B == 1'b1 && CI == 1'b1)
       (A *> S) = (tpllh$A$S$B_EQ_1_AN_CI_EQ_1, tphhl$A$S$B_EQ_1_AN_CI_EQ_1);
     if (B == 1'b1 && CI == 1'b0)
       (A *> S) = (tphlh$A$S$B_EQ_1_AN_CI_EQ_0, tplhl$A$S$B_EQ_1_AN_CI_EQ_0);
     if (B == 1'b0 && CI == 1'b1)
       (A *> S) = (tphlh$A$S$B_EQ_0_AN_CI_EQ_1, tplhl$A$S$B_EQ_0_AN_CI_EQ_1);
     if (B == 1'b0 && CI == 1'b0)
       (A *> S) = (tpllh$A$S$B_EQ_0_AN_CI_EQ_0, tphhl$A$S$B_EQ_0_AN_CI_EQ_0);
     ifnone
       (A *> S) = (tpllh$A$S,tplhl$A$S);

     if (B == 1'b1 && CI == 1'b0)
       (A *> CO) = (tpllh$A$CO$B_EQ_1_AN_CI_EQ_0, tphhl$A$CO$B_EQ_1_AN_CI_EQ_0);
     if (B == 1'b0 && CI == 1'b1)
       (A *> CO) = (tpllh$A$CO$B_EQ_0_AN_CI_EQ_1, tphhl$A$CO$B_EQ_0_AN_CI_EQ_1);
     ifnone
       (A *> CO) = (tpllh$A$CO,tphhl$A$CO);*/
 // path delays
      (posedge A => (S +: S)) = (1.0, 1.0);
      (negedge A => (S -: S)) = (1.0, 1.0);
      if (B == 1'b1 && CI == 1'b0) (A +=> CO) = (1.0, 1.0);
      if (B == 1'b0 && CI == 1'b1) (A +=> CO) = (1.0, 1.0);
 
      if (B == 1'b1 && CI == 1'b1) (A +=> S) = (1.0, 1.0);
      if (B == 1'b0 && CI == 1'b0) (A +=> S) = (1.0, 1.0);
      if (B == 1'b1 && CI == 1'b0) (A -=> S) = (1.0, 1.0);
      if (B == 1'b0 && CI == 1'b1) (A -=> S) = (1.0, 1.0);

   

      (posedge B => (S +: S)) = (1.0, 1.0);
      (negedge B => (S -: S)) = (1.0, 1.0);
      if (A == 1'b1 && CI == 1'b0) (B +=> CO) = (1.0, 1.0);
      if (A == 1'b0 && CI == 1'b1) (B +=> CO) = (1.0, 1.0);
  
      if (A == 1'b1 && CI == 1'b1) (B +=> S) = (1.0, 1.0);
      if (A == 1'b0 && CI == 1'b0) (B +=> S) = (1.0, 1.0);
      if (A == 1'b0 && CI == 1'b1) (B -=> S) = (1.0, 1.0);
      if (A == 1'b1 && CI == 1'b0) (B -=> S) = (1.0, 1.0);
   

      (posedge CI => (S +: S)) = (1.0, 1.0);
      (negedge CI => (S -: S)) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0) (CI +=> CO) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1) (CI +=> CO) = (1.0, 1.0);

      if (A == 1'b1 && B == 1'b1) (CI +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b0) (CI +=> S) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0) (CI -=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1) (CI -=> S) = (1.0, 1.0);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_FA01D2 (CO, S, A, B, CI);
input  A ;
input  B ;
input  CI ;
output CO ;
output S ;

   and (I0_out, A, B);
   and (I1_out, B, CI);
   and (I3_out, CI, A);
   or  (CO, I0_out, I1_out, I3_out);
   xor (I5_out, A, B);
   xor (S, I5_out, CI);

   specify
     // delay parameters
  /*   specparam
       tpllh$A$S = 1.0,
       tplhl$A$S = 1.0,
       tphlh$A$S = 1.0,
       tphhl$A$S = 1.0,
       tpllh$A$CO = 1.0,
       tphhl$A$CO = 1.0,
       tpllh$B$S = 1.0,
       tplhl$B$S = 1.0,
       tphlh$B$S = 1.0,
       tphhl$B$S = 1.0,
       tpllh$B$CO = 1.0,
       tphhl$B$CO = 1.0,
       tpllh$CI$S = 1.0,
       tplhl$CI$S = 1.0,
       tphlh$CI$S = 1.0,
       tphhl$CI$S = 1.0,
       tpllh$CI$CO = 1.0,
       tphhl$CI$CO = 1.0,
       tpllh$A$S$B_EQ_1_AN_CI_EQ_1 = 1.0,
       tphhl$A$S$B_EQ_1_AN_CI_EQ_1 = 1.0,
       tpllh$A$S$B_EQ_0_AN_CI_EQ_0 = 1.0,
       tphhl$A$S$B_EQ_0_AN_CI_EQ_0 = 1.0,
       tplhl$A$S$B_EQ_1_AN_CI_EQ_0 = 1.0,
       tphlh$A$S$B_EQ_1_AN_CI_EQ_0 = 1.0,
       tplhl$A$S$B_EQ_0_AN_CI_EQ_1 = 1.0,
       tphlh$A$S$B_EQ_0_AN_CI_EQ_1 = 1.0,
       tpllh$A$CO$B_EQ_1_AN_CI_EQ_0 = 1.0,
       tphhl$A$CO$B_EQ_1_AN_CI_EQ_0 = 1.0,
       tpllh$A$CO$B_EQ_0_AN_CI_EQ_1 = 1.0,
       tphhl$A$CO$B_EQ_0_AN_CI_EQ_1 = 1.0,
       tpllh$B$S$A_EQ_1_AN_CI_EQ_1 = 1.0,
       tphhl$B$S$A_EQ_1_AN_CI_EQ_1 = 1.0,
       tpllh$B$S$A_EQ_0_AN_CI_EQ_0 = 1.0,
       tphhl$B$S$A_EQ_0_AN_CI_EQ_0 = 1.0,
       tplhl$B$S$A_EQ_0_AN_CI_EQ_1 = 1.0,
       tphlh$B$S$A_EQ_0_AN_CI_EQ_1 = 1.0,
       tplhl$B$S$A_EQ_1_AN_CI_EQ_0 = 1.0,
       tphlh$B$S$A_EQ_1_AN_CI_EQ_0 = 1.0,
       tpllh$B$CO$A_EQ_1_AN_CI_EQ_0 = 1.0,
       tphhl$B$CO$A_EQ_1_AN_CI_EQ_0 = 1.0,
       tpllh$B$CO$A_EQ_0_AN_CI_EQ_1 = 1.0,
       tphhl$B$CO$A_EQ_0_AN_CI_EQ_1 = 1.0,
       tpllh$CI$S$A_EQ_1_AN_B_EQ_1 = 1.0,
       tphhl$CI$S$A_EQ_1_AN_B_EQ_1 = 1.0,
       tpllh$CI$S$A_EQ_0_AN_B_EQ_0 = 1.0,
       tphhl$CI$S$A_EQ_0_AN_B_EQ_0 = 1.0,
       tplhl$CI$S$A_EQ_1_AN_B_EQ_0 = 1.0,
       tphlh$CI$S$A_EQ_1_AN_B_EQ_0 = 1.0,
       tplhl$CI$S$A_EQ_0_AN_B_EQ_1 = 1.0,
       tphlh$CI$S$A_EQ_0_AN_B_EQ_1 = 1.0,
       tpllh$CI$CO$A_EQ_1_AN_B_EQ_0 = 1.0,
       tphhl$CI$CO$A_EQ_1_AN_B_EQ_0 = 1.0,
       tpllh$CI$CO$A_EQ_0_AN_B_EQ_1 = 1.0,
       tphhl$CI$CO$A_EQ_0_AN_B_EQ_1 = 1.0;

     // path delays
     if (A == 1'b1 && B == 1'b1)
       (CI *> S) = (tpllh$CI$S$A_EQ_1_AN_B_EQ_1, tphhl$CI$S$A_EQ_1_AN_B_EQ_1);
     if (A == 1'b1 && B == 1'b0)
       (CI *> S) = (tphlh$CI$S$A_EQ_1_AN_B_EQ_0, tplhl$CI$S$A_EQ_1_AN_B_EQ_0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> S) = (tphlh$CI$S$A_EQ_0_AN_B_EQ_1, tplhl$CI$S$A_EQ_0_AN_B_EQ_1);
     if (A == 1'b0 && B == 1'b0)
       (CI *> S) = (tpllh$CI$S$A_EQ_0_AN_B_EQ_0, tphhl$CI$S$A_EQ_0_AN_B_EQ_0);
     ifnone
       (CI *> S) = (tpllh$CI$S,tplhl$CI$S);

     if (A == 1'b1 && B == 1'b0)
       (CI *> CO) = (tpllh$CI$CO$A_EQ_1_AN_B_EQ_0, tphhl$CI$CO$A_EQ_1_AN_B_EQ_0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> CO) = (tpllh$CI$CO$A_EQ_0_AN_B_EQ_1, tphhl$CI$CO$A_EQ_0_AN_B_EQ_1);
     ifnone
       (CI *> CO) = (tpllh$CI$CO,tphhl$CI$CO);

     if (A == 1'b1 && CI == 1'b1)
       (B *> S) = (tpllh$B$S$A_EQ_1_AN_CI_EQ_1, tphhl$B$S$A_EQ_1_AN_CI_EQ_1);
     if (A == 1'b1 && CI == 1'b0)
       (B *> S) = (tphlh$B$S$A_EQ_1_AN_CI_EQ_0, tplhl$B$S$A_EQ_1_AN_CI_EQ_0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> S) = (tphlh$B$S$A_EQ_0_AN_CI_EQ_1, tplhl$B$S$A_EQ_0_AN_CI_EQ_1);
     if (A == 1'b0 && CI == 1'b0)
       (B *> S) = (tpllh$B$S$A_EQ_0_AN_CI_EQ_0, tphhl$B$S$A_EQ_0_AN_CI_EQ_0);
     ifnone
       (B *> S) = (tpllh$B$S,tplhl$B$S);

     if (A == 1'b1 && CI == 1'b0)
       (B *> CO) = (tpllh$B$CO$A_EQ_1_AN_CI_EQ_0, tphhl$B$CO$A_EQ_1_AN_CI_EQ_0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> CO) = (tpllh$B$CO$A_EQ_0_AN_CI_EQ_1, tphhl$B$CO$A_EQ_0_AN_CI_EQ_1);
     ifnone
       (B *> CO) = (tpllh$B$CO,tphhl$B$CO);

     if (B == 1'b1 && CI == 1'b1)
       (A *> S) = (tpllh$A$S$B_EQ_1_AN_CI_EQ_1, tphhl$A$S$B_EQ_1_AN_CI_EQ_1);
     if (B == 1'b1 && CI == 1'b0)
       (A *> S) = (tphlh$A$S$B_EQ_1_AN_CI_EQ_0, tplhl$A$S$B_EQ_1_AN_CI_EQ_0);
     if (B == 1'b0 && CI == 1'b1)
       (A *> S) = (tphlh$A$S$B_EQ_0_AN_CI_EQ_1, tplhl$A$S$B_EQ_0_AN_CI_EQ_1);
     if (B == 1'b0 && CI == 1'b0)
       (A *> S) = (tpllh$A$S$B_EQ_0_AN_CI_EQ_0, tphhl$A$S$B_EQ_0_AN_CI_EQ_0);
     ifnone
       (A *> S) = (tpllh$A$S,tplhl$A$S);

     if (B == 1'b1 && CI == 1'b0)
       (A *> CO) = (tpllh$A$CO$B_EQ_1_AN_CI_EQ_0, tphhl$A$CO$B_EQ_1_AN_CI_EQ_0);
     if (B == 1'b0 && CI == 1'b1)
       (A *> CO) = (tpllh$A$CO$B_EQ_0_AN_CI_EQ_1, tphhl$A$CO$B_EQ_0_AN_CI_EQ_1);
     ifnone
       (A *> CO) = (tpllh$A$CO,tphhl$A$CO);*/

 // path delays
      (posedge A => (S +: S)) = (1.0, 1.0);
      (negedge A => (S -: S)) = (1.0, 1.0);
      if (B == 1'b1 && CI == 1'b0) (A +=> CO) = (1.0, 1.0);
      if (B == 1'b0 && CI == 1'b1) (A +=> CO) = (1.0, 1.0);
 
      if (B == 1'b1 && CI == 1'b1) (A +=> S) = (1.0, 1.0);
      if (B == 1'b0 && CI == 1'b0) (A +=> S) = (1.0, 1.0);
      if (B == 1'b1 && CI == 1'b0) (A -=> S) = (1.0, 1.0);
      if (B == 1'b0 && CI == 1'b1) (A -=> S) = (1.0, 1.0);

   

      (posedge B => (S +: S)) = (1.0, 1.0);
      (negedge B => (S -: S)) = (1.0, 1.0);
      if (A == 1'b1 && CI == 1'b0) (B +=> CO) = (1.0, 1.0);
      if (A == 1'b0 && CI == 1'b1) (B +=> CO) = (1.0, 1.0);
  
      if (A == 1'b1 && CI == 1'b1) (B +=> S) = (1.0, 1.0);
      if (A == 1'b0 && CI == 1'b0) (B +=> S) = (1.0, 1.0);
      if (A == 1'b0 && CI == 1'b1) (B -=> S) = (1.0, 1.0);
      if (A == 1'b1 && CI == 1'b0) (B -=> S) = (1.0, 1.0);
   

      (posedge CI => (S +: S)) = (1.0, 1.0);
      (negedge CI => (S -: S)) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0) (CI +=> CO) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1) (CI +=> CO) = (1.0, 1.0);

      if (A == 1'b1 && B == 1'b1) (CI +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b0) (CI +=> S) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0) (CI -=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1) (CI -=> S) = (1.0, 1.0);



   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_FA01D4 (CO, S, A, B, CI);
input  A ;
input  B ;
input  CI ;
output CO ;
output S ;

   and (I0_out, A, B);
   and (I1_out, B, CI);
   and (I3_out, CI, A);
   or  (CO, I0_out, I1_out, I3_out);
   xor (I5_out, A, B);
   xor (S, I5_out, CI);

   specify
     // delay parameters
   /*  specparam
       tpllh$A$S = 1.0,
       tplhl$A$S = 1.0,
       tphlh$A$S = 1.0,
       tphhl$A$S = 1.0,
       tpllh$A$CO = 1.0,
       tphhl$A$CO = 1.0,
       tpllh$B$S = 1.0,
       tplhl$B$S = 1.0,
       tphlh$B$S = 1.0,
       tphhl$B$S = 1.0,
       tpllh$B$CO = 1.0,
       tphhl$B$CO = 1.0,
       tpllh$CI$S = 1.0,
       tplhl$CI$S = 1.0,
       tphlh$CI$S = 1.0,
       tphhl$CI$S = 1.0,
       tpllh$CI$CO = 1.0,
       tphhl$CI$CO = 1.0,
       tpllh$A$S$B_EQ_1_AN_CI_EQ_1 = 1.0,
       tphhl$A$S$B_EQ_1_AN_CI_EQ_1 = 1.0,
       tpllh$A$S$B_EQ_0_AN_CI_EQ_0 = 1.0,
       tphhl$A$S$B_EQ_0_AN_CI_EQ_0 = 1.0,
       tplhl$A$S$B_EQ_1_AN_CI_EQ_0 = 1.0,
       tphlh$A$S$B_EQ_1_AN_CI_EQ_0 = 1.0,
       tplhl$A$S$B_EQ_0_AN_CI_EQ_1 = 1.0,
       tphlh$A$S$B_EQ_0_AN_CI_EQ_1 = 1.0,
       tpllh$A$CO$B_EQ_1_AN_CI_EQ_0 = 1.0,
       tphhl$A$CO$B_EQ_1_AN_CI_EQ_0 = 1.0,
       tpllh$A$CO$B_EQ_0_AN_CI_EQ_1 = 1.0,
       tphhl$A$CO$B_EQ_0_AN_CI_EQ_1 = 1.0,
       tpllh$B$S$A_EQ_1_AN_CI_EQ_1 = 1.0,
       tphhl$B$S$A_EQ_1_AN_CI_EQ_1 = 1.0,
       tpllh$B$S$A_EQ_0_AN_CI_EQ_0 = 1.0,
       tphhl$B$S$A_EQ_0_AN_CI_EQ_0 = 1.0,
       tplhl$B$S$A_EQ_0_AN_CI_EQ_1 = 1.0,
       tphlh$B$S$A_EQ_0_AN_CI_EQ_1 = 1.0,
       tplhl$B$S$A_EQ_1_AN_CI_EQ_0 = 1.0,
       tphlh$B$S$A_EQ_1_AN_CI_EQ_0 = 1.0,
       tpllh$B$CO$A_EQ_1_AN_CI_EQ_0 = 1.0,
       tphhl$B$CO$A_EQ_1_AN_CI_EQ_0 = 1.0,
       tpllh$B$CO$A_EQ_0_AN_CI_EQ_1 = 1.0,
       tphhl$B$CO$A_EQ_0_AN_CI_EQ_1 = 1.0,
       tpllh$CI$S$A_EQ_1_AN_B_EQ_1 = 1.0,
       tphhl$CI$S$A_EQ_1_AN_B_EQ_1 = 1.0,
       tpllh$CI$S$A_EQ_0_AN_B_EQ_0 = 1.0,
       tphhl$CI$S$A_EQ_0_AN_B_EQ_0 = 1.0,
       tplhl$CI$S$A_EQ_1_AN_B_EQ_0 = 1.0,
       tphlh$CI$S$A_EQ_1_AN_B_EQ_0 = 1.0,
       tplhl$CI$S$A_EQ_0_AN_B_EQ_1 = 1.0,
       tphlh$CI$S$A_EQ_0_AN_B_EQ_1 = 1.0,
       tpllh$CI$CO$A_EQ_1_AN_B_EQ_0 = 1.0,
       tphhl$CI$CO$A_EQ_1_AN_B_EQ_0 = 1.0,
       tpllh$CI$CO$A_EQ_0_AN_B_EQ_1 = 1.0,
       tphhl$CI$CO$A_EQ_0_AN_B_EQ_1 = 1.0;

     // path delays
     if (A == 1'b1 && B == 1'b1)
       (CI *> S) = (tpllh$CI$S$A_EQ_1_AN_B_EQ_1, tphhl$CI$S$A_EQ_1_AN_B_EQ_1);
     if (A == 1'b1 && B == 1'b0)
       (CI *> S) = (tphlh$CI$S$A_EQ_1_AN_B_EQ_0, tplhl$CI$S$A_EQ_1_AN_B_EQ_0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> S) = (tphlh$CI$S$A_EQ_0_AN_B_EQ_1, tplhl$CI$S$A_EQ_0_AN_B_EQ_1);
     if (A == 1'b0 && B == 1'b0)
       (CI *> S) = (tpllh$CI$S$A_EQ_0_AN_B_EQ_0, tphhl$CI$S$A_EQ_0_AN_B_EQ_0);
     ifnone
       (CI *> S) = (tpllh$CI$S,tplhl$CI$S);

     if (A == 1'b1 && B == 1'b0)
       (CI *> CO) = (tpllh$CI$CO$A_EQ_1_AN_B_EQ_0, tphhl$CI$CO$A_EQ_1_AN_B_EQ_0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> CO) = (tpllh$CI$CO$A_EQ_0_AN_B_EQ_1, tphhl$CI$CO$A_EQ_0_AN_B_EQ_1);
     ifnone
       (CI *> CO) = (tpllh$CI$CO,tphhl$CI$CO);

     if (A == 1'b1 && CI == 1'b1)
       (B *> S) = (tpllh$B$S$A_EQ_1_AN_CI_EQ_1, tphhl$B$S$A_EQ_1_AN_CI_EQ_1);
     if (A == 1'b1 && CI == 1'b0)
       (B *> S) = (tphlh$B$S$A_EQ_1_AN_CI_EQ_0, tplhl$B$S$A_EQ_1_AN_CI_EQ_0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> S) = (tphlh$B$S$A_EQ_0_AN_CI_EQ_1, tplhl$B$S$A_EQ_0_AN_CI_EQ_1);
     if (A == 1'b0 && CI == 1'b0)
       (B *> S) = (tpllh$B$S$A_EQ_0_AN_CI_EQ_0, tphhl$B$S$A_EQ_0_AN_CI_EQ_0);
     ifnone
       (B *> S) = (tpllh$B$S,tplhl$B$S);

     if (A == 1'b1 && CI == 1'b0)
       (B *> CO) = (tpllh$B$CO$A_EQ_1_AN_CI_EQ_0, tphhl$B$CO$A_EQ_1_AN_CI_EQ_0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> CO) = (tpllh$B$CO$A_EQ_0_AN_CI_EQ_1, tphhl$B$CO$A_EQ_0_AN_CI_EQ_1);
     ifnone
       (B *> CO) = (tpllh$B$CO,tphhl$B$CO);

     if (B == 1'b1 && CI == 1'b1)
       (A *> S) = (tpllh$A$S$B_EQ_1_AN_CI_EQ_1, tphhl$A$S$B_EQ_1_AN_CI_EQ_1);
     if (B == 1'b1 && CI == 1'b0)
       (A *> S) = (tphlh$A$S$B_EQ_1_AN_CI_EQ_0, tplhl$A$S$B_EQ_1_AN_CI_EQ_0);
     if (B == 1'b0 && CI == 1'b1)
       (A *> S) = (tphlh$A$S$B_EQ_0_AN_CI_EQ_1, tplhl$A$S$B_EQ_0_AN_CI_EQ_1);
     if (B == 1'b0 && CI == 1'b0)
       (A *> S) = (tpllh$A$S$B_EQ_0_AN_CI_EQ_0, tphhl$A$S$B_EQ_0_AN_CI_EQ_0);
     ifnone
       (A *> S) = (tpllh$A$S,tplhl$A$S);

     if (B == 1'b1 && CI == 1'b0)
       (A *> CO) = (tpllh$A$CO$B_EQ_1_AN_CI_EQ_0, tphhl$A$CO$B_EQ_1_AN_CI_EQ_0);
     if (B == 1'b0 && CI == 1'b1)
       (A *> CO) = (tpllh$A$CO$B_EQ_0_AN_CI_EQ_1, tphhl$A$CO$B_EQ_0_AN_CI_EQ_1);
     ifnone
       (A *> CO) = (tpllh$A$CO,tphhl$A$CO);*/

// path delays
      (posedge A => (S +: S)) = (1.0, 1.0);
      (negedge A => (S -: S)) = (1.0, 1.0);
      if (B == 1'b1 && CI == 1'b0) (A +=> CO) = (1.0, 1.0);
      if (B == 1'b0 && CI == 1'b1) (A +=> CO) = (1.0, 1.0);
 
      if (B == 1'b1 && CI == 1'b1) (A +=> S) = (1.0, 1.0);
      if (B == 1'b0 && CI == 1'b0) (A +=> S) = (1.0, 1.0);
      if (B == 1'b1 && CI == 1'b0) (A -=> S) = (1.0, 1.0);
      if (B == 1'b0 && CI == 1'b1) (A -=> S) = (1.0, 1.0);

   

      (posedge B => (S +: S)) = (1.0, 1.0);
      (negedge B => (S -: S)) = (1.0, 1.0);
      if (A == 1'b1 && CI == 1'b0) (B +=> CO) = (1.0, 1.0);
      if (A == 1'b0 && CI == 1'b1) (B +=> CO) = (1.0, 1.0);
  
      if (A == 1'b1 && CI == 1'b1) (B +=> S) = (1.0, 1.0);
      if (A == 1'b0 && CI == 1'b0) (B +=> S) = (1.0, 1.0);
      if (A == 1'b0 && CI == 1'b1) (B -=> S) = (1.0, 1.0);
      if (A == 1'b1 && CI == 1'b0) (B -=> S) = (1.0, 1.0);
   

      (posedge CI => (S +: S)) = (1.0, 1.0);
      (negedge CI => (S -: S)) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0) (CI +=> CO) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1) (CI +=> CO) = (1.0, 1.0);

      if (A == 1'b1 && B == 1'b1) (CI +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b0) (CI +=> S) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0) (CI -=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1) (CI -=> S) = (1.0, 1.0);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_FA02D1 (NCO, S, A, B, CI);
input  A ;
input  B ;
input  CI ;
output NCO ;
output S ;

   and (I0_out, A, B);
   and (I1_out, B, CI);
   and (I3_out, CI, A);
   or  (I4_out, I0_out, I1_out, I3_out);
   not (NCO, I4_out);
   xor (I6_out, A, B);
   xor (S, I6_out, CI);

   specify
     // delay parameters
    /*  specparam
       tpllh$A$S = 1.0,
       tplhl$A$S = 1.0,
       tphlh$A$S = 1.0,
       tphhl$A$S = 1.0,
       tplhl$A$NCO = 1.0,
       tphlh$A$NCO = 1.0,
       tpllh$B$S = 1.0,
       tplhl$B$S = 1.0,
       tphlh$B$S = 1.0,
       tphhl$B$S = 1.0,
       tplhl$B$NCO = 1.0,
       tphlh$B$NCO = 1.0,
       tpllh$CI$S = 1.0,
       tplhl$CI$S = 1.0,
       tphlh$CI$S = 1.0,
       tphhl$CI$S = 1.0,
       tplhl$CI$NCO = 1.0,
       tphlh$CI$NCO = 1.0,
       tpllh$A$S$B_EQ_1_AN_CI_EQ_1 = 1.0,
       tphhl$A$S$B_EQ_1_AN_CI_EQ_1 = 1.0,
       tpllh$A$S$B_EQ_0_AN_CI_EQ_0 = 1.0,
       tphhl$A$S$B_EQ_0_AN_CI_EQ_0 = 1.0,
       tplhl$A$S$B_EQ_1_AN_CI_EQ_0 = 1.0,
       tphlh$A$S$B_EQ_1_AN_CI_EQ_0 = 1.0,
       tplhl$A$S$B_EQ_0_AN_CI_EQ_1 = 1.0,
       tphlh$A$S$B_EQ_0_AN_CI_EQ_1 = 1.0,
       tplhl$A$NCO$B_EQ_1_AN_CI_EQ_0 = 1.0,
       tphlh$A$NCO$B_EQ_1_AN_CI_EQ_0 = 1.0,
       tplhl$A$NCO$B_EQ_0_AN_CI_EQ_1 = 1.0,
       tphlh$A$NCO$B_EQ_0_AN_CI_EQ_1 = 1.0,
       tpllh$B$S$A_EQ_1_AN_CI_EQ_1 = 1.0,
       tphhl$B$S$A_EQ_1_AN_CI_EQ_1 = 1.0,
       tpllh$B$S$A_EQ_0_AN_CI_EQ_0 = 1.0,
       tphhl$B$S$A_EQ_0_AN_CI_EQ_0 = 1.0,
       tplhl$B$S$A_EQ_1_AN_CI_EQ_0 = 1.0,
       tphlh$B$S$A_EQ_1_AN_CI_EQ_0 = 1.0,
       tplhl$B$S$A_EQ_0_AN_CI_EQ_1 = 1.0,
       tphlh$B$S$A_EQ_0_AN_CI_EQ_1 = 1.0,
       tplhl$B$NCO$A_EQ_1_AN_CI_EQ_0 = 1.0,
       tphlh$B$NCO$A_EQ_1_AN_CI_EQ_0 = 1.0,
       tplhl$B$NCO$A_EQ_0_AN_CI_EQ_1 = 1.0,
       tphlh$B$NCO$A_EQ_0_AN_CI_EQ_1 = 1.0,
       tpllh$CI$S$A_EQ_1_AN_B_EQ_1 = 1.0,
       tphhl$CI$S$A_EQ_1_AN_B_EQ_1 = 1.0,
       tpllh$CI$S$A_EQ_0_AN_B_EQ_0 = 1.0,
       tphhl$CI$S$A_EQ_0_AN_B_EQ_0 = 1.0,
       tplhl$CI$S$A_EQ_1_AN_B_EQ_0 = 1.0,
       tphlh$CI$S$A_EQ_1_AN_B_EQ_0 = 1.0,
       tplhl$CI$S$A_EQ_0_AN_B_EQ_1 = 1.0,
       tphlh$CI$S$A_EQ_0_AN_B_EQ_1 = 1.0,
       tplhl$CI$NCO$A_EQ_1_AN_B_EQ_0 = 1.0,
       tphlh$CI$NCO$A_EQ_1_AN_B_EQ_0 = 1.0,
       tplhl$CI$NCO$A_EQ_0_AN_B_EQ_1 = 1.0,
       tphlh$CI$NCO$A_EQ_0_AN_B_EQ_1 = 1.0;

     // path delays
    if (A == 1'b1 && B == 1'b1)
       (CI *> S) = (tpllh$CI$S$A_EQ_1_AN_B_EQ_1, tphhl$CI$S$A_EQ_1_AN_B_EQ_1);
     if (A == 1'b1 && B == 1'b0)
       (CI *> S) = (tphlh$CI$S$A_EQ_1_AN_B_EQ_0, tplhl$CI$S$A_EQ_1_AN_B_EQ_0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> S) = (tphlh$CI$S$A_EQ_0_AN_B_EQ_1, tplhl$CI$S$A_EQ_0_AN_B_EQ_1);
     if (A == 1'b0 && B == 1'b0)
       (CI *> S) = (tpllh$CI$S$A_EQ_0_AN_B_EQ_0, tphhl$CI$S$A_EQ_0_AN_B_EQ_0);
     ifnone
       (CI *> S) = (tpllh$CI$S,tplhl$CI$S);

     if (A == 1'b1 && B == 1'b0)
       (CI *> NCO) = (tphlh$CI$NCO$A_EQ_1_AN_B_EQ_0, tplhl$CI$NCO$A_EQ_1_AN_B_EQ_0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> NCO) = (tphlh$CI$NCO$A_EQ_0_AN_B_EQ_1, tplhl$CI$NCO$A_EQ_0_AN_B_EQ_1);
     ifnone
       (CI *> NCO) = (tphlh$CI$NCO,tplhl$CI$NCO);

     if (A == 1'b1 && CI == 1'b1)
       (B *> S) = (tpllh$B$S$A_EQ_1_AN_CI_EQ_1, tphhl$B$S$A_EQ_1_AN_CI_EQ_1);
     if (A == 1'b1 && CI == 1'b0)
       (B *> S) = (tphlh$B$S$A_EQ_1_AN_CI_EQ_0, tplhl$B$S$A_EQ_1_AN_CI_EQ_0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> S) = (tphlh$B$S$A_EQ_0_AN_CI_EQ_1, tplhl$B$S$A_EQ_0_AN_CI_EQ_1);
     if (A == 1'b0 && CI == 1'b0)
       (B *> S) = (tpllh$B$S$A_EQ_0_AN_CI_EQ_0, tphhl$B$S$A_EQ_0_AN_CI_EQ_0);
     ifnone
       (B *> S) = (tpllh$B$S,tplhl$B$S);

     if (A == 1'b1 && CI == 1'b0)
       (B *> NCO) = (tphlh$B$NCO$A_EQ_1_AN_CI_EQ_0, tplhl$B$NCO$A_EQ_1_AN_CI_EQ_0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> NCO) = (tphlh$B$NCO$A_EQ_0_AN_CI_EQ_1, tplhl$B$NCO$A_EQ_0_AN_CI_EQ_1);
     ifnone
       (B *> NCO) = (tphlh$B$NCO,tplhl$B$NCO);

     if (B == 1'b1 && CI == 1'b1)
       (A *> S) = (tpllh$A$S$B_EQ_1_AN_CI_EQ_1, tphhl$A$S$B_EQ_1_AN_CI_EQ_1);
     if (B == 1'b1 && CI == 1'b0)
       (A *> S) = (tphlh$A$S$B_EQ_1_AN_CI_EQ_0, tplhl$A$S$B_EQ_1_AN_CI_EQ_0);
     if (B == 1'b0 && CI == 1'b1)
       (A *> S) = (tphlh$A$S$B_EQ_0_AN_CI_EQ_1, tplhl$A$S$B_EQ_0_AN_CI_EQ_1);
     if (B == 1'b0 && CI == 1'b0)
       (A *> S) = (tpllh$A$S$B_EQ_0_AN_CI_EQ_0, tphhl$A$S$B_EQ_0_AN_CI_EQ_0);
     ifnone
       (A *> S) = (tpllh$A$S,tplhl$A$S);

     if (B == 1'b1 && CI == 1'b0)
       (A *> NCO) = (tphlh$A$NCO$B_EQ_1_AN_CI_EQ_0, tplhl$A$NCO$B_EQ_1_AN_CI_EQ_0);
     if (B == 1'b0 && CI == 1'b1)
       (A *> NCO) = (tphlh$A$NCO$B_EQ_0_AN_CI_EQ_1, tplhl$A$NCO$B_EQ_0_AN_CI_EQ_1);
     ifnone
       (A *> NCO) = (tphlh$A$NCO,tplhl$A$NCO);*/


// path delays
      (posedge A => (NCO +: NCO)) = (1.0, 1.0);
      (negedge A => (NCO -: NCO)) = (1.0, 1.0);
      if (B == 1'b1 && CI == 1'b0) (A -=> NCO) = (1.0, 1.0);
      if (B == 1'b0 && CI == 1'b1) (A -=> NCO) = (1.0, 1.0);
 
      if (B == 1'b1 && CI == 1'b1) (A +=> S) = (1.0, 1.0);
      if (B == 1'b0 && CI == 1'b0) (A +=> S) = (1.0, 1.0);
      if (B == 1'b1 && CI == 1'b0) (A -=> S) = (1.0, 1.0);
      if (B == 1'b0 && CI == 1'b1) (A -=> S) = (1.0, 1.0);

   

      (posedge B => (S +: S)) = (1.0, 1.0);
      (negedge B => (S -: S)) = (1.0, 1.0);
      if (A == 1'b1 && CI == 1'b0) (B -=> NCO) = (1.0, 1.0);
      if (A == 1'b0 && CI == 1'b1) (B -=> NCO) = (1.0, 1.0);
  
      if (A == 1'b1 && CI == 1'b1) (B +=> S) = (1.0, 1.0);
      if (A == 1'b0 && CI == 1'b0) (B +=> S) = (1.0, 1.0);
      if (A == 1'b0 && CI == 1'b1) (B -=> S) = (1.0, 1.0);
      if (A == 1'b1 && CI == 1'b0) (B -=> S) = (1.0, 1.0);
   

      (posedge CI => (S +: S)) = (1.0, 1.0);
      (negedge CI => (S -: S)) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0) (CI +=> NCO) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1) (CI +=> NCO) = (1.0, 1.0);

      if (A == 1'b1 && B == 1'b1) (CI +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b0) (CI +=> S) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0) (CI -=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1) (CI -=> S) = (1.0, 1.0);






   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_FA02D2 (NCO, S, A, B, CI);
input  A ;
input  B ;
input  CI ;
output NCO ;
output S ;

   and (I0_out, A, B);
   and (I1_out, B, CI);
   and (I3_out, CI, A);
   or  (I4_out, I0_out, I1_out, I3_out);
   not (NCO, I4_out);
   xor (I6_out, A, B);
   xor (S, I6_out, CI);

   specify
     // delay parameters
  /*   specparam
       tpllh$A$S = 1.0,
       tplhl$A$S = 1.0,
       tphlh$A$S = 1.0,
       tphhl$A$S = 1.0,
       tplhl$A$NCO = 1.0,
       tphlh$A$NCO = 1.0,
       tpllh$B$S = 1.0,
       tplhl$B$S = 1.0,
       tphlh$B$S = 1.0,
       tphhl$B$S = 1.0,
       tplhl$B$NCO = 1.0,
       tphlh$B$NCO = 1.0,
       tpllh$CI$S = 1.0,
       tplhl$CI$S = 1.0,
       tphlh$CI$S = 1.0,
       tphhl$CI$S = 1.0,
       tplhl$CI$NCO = 1.0,
       tphlh$CI$NCO = 1.0,
       tpllh$A$S$B_EQ_1_AN_CI_EQ_1 = 1.0,
       tphhl$A$S$B_EQ_1_AN_CI_EQ_1 = 1.0,
       tpllh$A$S$B_EQ_0_AN_CI_EQ_0 = 1.0,
       tphhl$A$S$B_EQ_0_AN_CI_EQ_0 = 1.0,
       tplhl$A$S$B_EQ_1_AN_CI_EQ_0 = 1.0,
       tphlh$A$S$B_EQ_1_AN_CI_EQ_0 = 1.0,
       tplhl$A$S$B_EQ_0_AN_CI_EQ_1 = 1.0,
       tphlh$A$S$B_EQ_0_AN_CI_EQ_1 = 1.0,
       tplhl$A$NCO$B_EQ_1_AN_CI_EQ_0 = 1.0,
       tphlh$A$NCO$B_EQ_1_AN_CI_EQ_0 = 1.0,
       tplhl$A$NCO$B_EQ_0_AN_CI_EQ_1 = 1.0,
       tphlh$A$NCO$B_EQ_0_AN_CI_EQ_1 = 1.0,
       tpllh$B$S$A_EQ_1_AN_CI_EQ_1 = 1.0,
       tphhl$B$S$A_EQ_1_AN_CI_EQ_1 = 1.0,
       tpllh$B$S$A_EQ_0_AN_CI_EQ_0 = 1.0,
       tphhl$B$S$A_EQ_0_AN_CI_EQ_0 = 1.0,
       tplhl$B$S$A_EQ_1_AN_CI_EQ_0 = 1.0,
       tphlh$B$S$A_EQ_1_AN_CI_EQ_0 = 1.0,
       tplhl$B$S$A_EQ_0_AN_CI_EQ_1 = 1.0,
       tphlh$B$S$A_EQ_0_AN_CI_EQ_1 = 1.0,
       tplhl$B$NCO$A_EQ_1_AN_CI_EQ_0 = 1.0,
       tphlh$B$NCO$A_EQ_1_AN_CI_EQ_0 = 1.0,
       tplhl$B$NCO$A_EQ_0_AN_CI_EQ_1 = 1.0,
       tphlh$B$NCO$A_EQ_0_AN_CI_EQ_1 = 1.0,
       tpllh$CI$S$A_EQ_1_AN_B_EQ_1 = 1.0,
       tphhl$CI$S$A_EQ_1_AN_B_EQ_1 = 1.0,
       tpllh$CI$S$A_EQ_0_AN_B_EQ_0 = 1.0,
       tphhl$CI$S$A_EQ_0_AN_B_EQ_0 = 1.0,
       tplhl$CI$S$A_EQ_1_AN_B_EQ_0 = 1.0,
       tphlh$CI$S$A_EQ_1_AN_B_EQ_0 = 1.0,
       tplhl$CI$S$A_EQ_0_AN_B_EQ_1 = 1.0,
       tphlh$CI$S$A_EQ_0_AN_B_EQ_1 = 1.0,
       tplhl$CI$NCO$A_EQ_1_AN_B_EQ_0 = 1.0,
       tphlh$CI$NCO$A_EQ_1_AN_B_EQ_0 = 1.0,
       tplhl$CI$NCO$A_EQ_0_AN_B_EQ_1 = 1.0,
       tphlh$CI$NCO$A_EQ_0_AN_B_EQ_1 = 1.0;

     // path delays
     if (A == 1'b1 && B == 1'b1)
       (CI *> S) = (tpllh$CI$S$A_EQ_1_AN_B_EQ_1, tphhl$CI$S$A_EQ_1_AN_B_EQ_1);
     if (A == 1'b1 && B == 1'b0)
       (CI *> S) = (tphlh$CI$S$A_EQ_1_AN_B_EQ_0, tplhl$CI$S$A_EQ_1_AN_B_EQ_0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> S) = (tphlh$CI$S$A_EQ_0_AN_B_EQ_1, tplhl$CI$S$A_EQ_0_AN_B_EQ_1);
     if (A == 1'b0 && B == 1'b0)
       (CI *> S) = (tpllh$CI$S$A_EQ_0_AN_B_EQ_0, tphhl$CI$S$A_EQ_0_AN_B_EQ_0);
     ifnone
       (CI *> S) = (tpllh$CI$S,tplhl$CI$S);

     if (A == 1'b1 && B == 1'b0)
       (CI *> NCO) = (tphlh$CI$NCO$A_EQ_1_AN_B_EQ_0, tplhl$CI$NCO$A_EQ_1_AN_B_EQ_0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> NCO) = (tphlh$CI$NCO$A_EQ_0_AN_B_EQ_1, tplhl$CI$NCO$A_EQ_0_AN_B_EQ_1);
     ifnone
       (CI *> NCO) = (tphlh$CI$NCO,tplhl$CI$NCO);

     if (A == 1'b1 && CI == 1'b1)
       (B *> S) = (tpllh$B$S$A_EQ_1_AN_CI_EQ_1, tphhl$B$S$A_EQ_1_AN_CI_EQ_1);
     if (A == 1'b1 && CI == 1'b0)
       (B *> S) = (tphlh$B$S$A_EQ_1_AN_CI_EQ_0, tplhl$B$S$A_EQ_1_AN_CI_EQ_0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> S) = (tphlh$B$S$A_EQ_0_AN_CI_EQ_1, tplhl$B$S$A_EQ_0_AN_CI_EQ_1);
     if (A == 1'b0 && CI == 1'b0)
       (B *> S) = (tpllh$B$S$A_EQ_0_AN_CI_EQ_0, tphhl$B$S$A_EQ_0_AN_CI_EQ_0);
     ifnone
       (B *> S) = (tpllh$B$S,tplhl$B$S);

     if (A == 1'b1 && CI == 1'b0)
       (B *> NCO) = (tphlh$B$NCO$A_EQ_1_AN_CI_EQ_0, tplhl$B$NCO$A_EQ_1_AN_CI_EQ_0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> NCO) = (tphlh$B$NCO$A_EQ_0_AN_CI_EQ_1, tplhl$B$NCO$A_EQ_0_AN_CI_EQ_1);
     ifnone
       (B *> NCO) = (tphlh$B$NCO,tplhl$B$NCO);

     if (B == 1'b1 && CI == 1'b1)
       (A *> S) = (tpllh$A$S$B_EQ_1_AN_CI_EQ_1, tphhl$A$S$B_EQ_1_AN_CI_EQ_1);
     if (B == 1'b1 && CI == 1'b0)
       (A *> S) = (tphlh$A$S$B_EQ_1_AN_CI_EQ_0, tplhl$A$S$B_EQ_1_AN_CI_EQ_0);
     if (B == 1'b0 && CI == 1'b1)
       (A *> S) = (tphlh$A$S$B_EQ_0_AN_CI_EQ_1, tplhl$A$S$B_EQ_0_AN_CI_EQ_1);
     if (B == 1'b0 && CI == 1'b0)
       (A *> S) = (tpllh$A$S$B_EQ_0_AN_CI_EQ_0, tphhl$A$S$B_EQ_0_AN_CI_EQ_0);
     ifnone
       (A *> S) = (tpllh$A$S,tplhl$A$S);

     if (B == 1'b1 && CI == 1'b0)
       (A *> NCO) = (tphlh$A$NCO$B_EQ_1_AN_CI_EQ_0, tplhl$A$NCO$B_EQ_1_AN_CI_EQ_0);
     if (B == 1'b0 && CI == 1'b1)
       (A *> NCO) = (tphlh$A$NCO$B_EQ_0_AN_CI_EQ_1, tplhl$A$NCO$B_EQ_0_AN_CI_EQ_1);
     ifnone
       (A *> NCO) = (tphlh$A$NCO,tplhl$A$NCO);*/

// path delays
      (posedge A => (NCO +: NCO)) = (1.0, 1.0);
      (negedge A => (NCO -: NCO)) = (1.0, 1.0);
      if (B == 1'b1 && CI == 1'b0) (A -=> NCO) = (1.0, 1.0);
      if (B == 1'b0 && CI == 1'b1) (A -=> NCO) = (1.0, 1.0);
 
      if (B == 1'b1 && CI == 1'b1) (A +=> S) = (1.0, 1.0);
      if (B == 1'b0 && CI == 1'b0) (A +=> S) = (1.0, 1.0);
      if (B == 1'b1 && CI == 1'b0) (A -=> S) = (1.0, 1.0);
      if (B == 1'b0 && CI == 1'b1) (A -=> S) = (1.0, 1.0);

   

      (posedge B => (S +: S)) = (1.0, 1.0);
      (negedge B => (S -: S)) = (1.0, 1.0);
      if (A == 1'b1 && CI == 1'b0) (B -=> NCO) = (1.0, 1.0);
      if (A == 1'b0 && CI == 1'b1) (B -=> NCO) = (1.0, 1.0);
  
      if (A == 1'b1 && CI == 1'b1) (B +=> S) = (1.0, 1.0);
      if (A == 1'b0 && CI == 1'b0) (B +=> S) = (1.0, 1.0);
      if (A == 1'b0 && CI == 1'b1) (B -=> S) = (1.0, 1.0);
      if (A == 1'b1 && CI == 1'b0) (B -=> S) = (1.0, 1.0);
   

      (posedge CI => (S +: S)) = (1.0, 1.0);
      (negedge CI => (S -: S)) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0) (CI +=> NCO) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1) (CI +=> NCO) = (1.0, 1.0);

      if (A == 1'b1 && B == 1'b1) (CI +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b0) (CI +=> S) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0) (CI -=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1) (CI -=> S) = (1.0, 1.0);


   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_FA02D4 (NCO, S, A, B, CI);
input  A ;
input  B ;
input  CI ;
output NCO ;
output S ;

   and (I0_out, A, B);
   and (I1_out, B, CI);
   and (I3_out, CI, A);
   or  (I4_out, I0_out, I1_out, I3_out);
   not (NCO, I4_out);
   xor (I6_out, A, B);
   xor (S, I6_out, CI);

   specify
     // delay parameters
  /*   specparam
       tpllh$A$S = 1.0,
       tplhl$A$S = 1.0,
       tphlh$A$S = 1.0,
       tphhl$A$S = 1.0,
       tplhl$A$NCO = 1.0,
       tphlh$A$NCO = 1.0,
       tpllh$B$S = 1.0,
       tplhl$B$S = 1.0,
       tphlh$B$S = 1.0,
       tphhl$B$S = 1.0,
       tplhl$B$NCO = 1.0,
       tphlh$B$NCO = 1.0,
       tpllh$CI$S = 1.0,
       tplhl$CI$S = 1.0,
       tphlh$CI$S = 1.0,
       tphhl$CI$S = 1.0,
       tplhl$CI$NCO = 1.0,
       tphlh$CI$NCO = 1.0,
       tpllh$A$S$B_EQ_1_AN_CI_EQ_1 = 1.0,
       tphhl$A$S$B_EQ_1_AN_CI_EQ_1 = 1.0,
       tpllh$A$S$B_EQ_0_AN_CI_EQ_0 = 1.0,
       tphhl$A$S$B_EQ_0_AN_CI_EQ_0 = 1.0,
       tplhl$A$S$B_EQ_1_AN_CI_EQ_0 = 1.0,
       tphlh$A$S$B_EQ_1_AN_CI_EQ_0 = 1.0,
       tplhl$A$S$B_EQ_0_AN_CI_EQ_1 = 1.0,
       tphlh$A$S$B_EQ_0_AN_CI_EQ_1 = 1.0,
       tplhl$A$NCO$B_EQ_1_AN_CI_EQ_0 = 1.0,
       tphlh$A$NCO$B_EQ_1_AN_CI_EQ_0 = 1.0,
       tplhl$A$NCO$B_EQ_0_AN_CI_EQ_1 = 1.0,
       tphlh$A$NCO$B_EQ_0_AN_CI_EQ_1 = 1.0,
       tpllh$B$S$A_EQ_1_AN_CI_EQ_1 = 1.0,
       tphhl$B$S$A_EQ_1_AN_CI_EQ_1 = 1.0,
       tpllh$B$S$A_EQ_0_AN_CI_EQ_0 = 1.0,
       tphhl$B$S$A_EQ_0_AN_CI_EQ_0 = 1.0,
       tplhl$B$S$A_EQ_1_AN_CI_EQ_0 = 1.0,
       tphlh$B$S$A_EQ_1_AN_CI_EQ_0 = 1.0,
       tplhl$B$S$A_EQ_0_AN_CI_EQ_1 = 1.0,
       tphlh$B$S$A_EQ_0_AN_CI_EQ_1 = 1.0,
       tplhl$B$NCO$A_EQ_1_AN_CI_EQ_0 = 1.0,
       tphlh$B$NCO$A_EQ_1_AN_CI_EQ_0 = 1.0,
       tplhl$B$NCO$A_EQ_0_AN_CI_EQ_1 = 1.0,
       tphlh$B$NCO$A_EQ_0_AN_CI_EQ_1 = 1.0,
       tpllh$CI$S$A_EQ_1_AN_B_EQ_1 = 1.0,
       tphhl$CI$S$A_EQ_1_AN_B_EQ_1 = 1.0,
       tpllh$CI$S$A_EQ_0_AN_B_EQ_0 = 1.0,
       tphhl$CI$S$A_EQ_0_AN_B_EQ_0 = 1.0,
       tplhl$CI$S$A_EQ_1_AN_B_EQ_0 = 1.0,
       tphlh$CI$S$A_EQ_1_AN_B_EQ_0 = 1.0,
       tplhl$CI$S$A_EQ_0_AN_B_EQ_1 = 1.0,
       tphlh$CI$S$A_EQ_0_AN_B_EQ_1 = 1.0,
       tplhl$CI$NCO$A_EQ_1_AN_B_EQ_0 = 1.0,
       tphlh$CI$NCO$A_EQ_1_AN_B_EQ_0 = 1.0,
       tplhl$CI$NCO$A_EQ_0_AN_B_EQ_1 = 1.0,
       tphlh$CI$NCO$A_EQ_0_AN_B_EQ_1 = 1.0;

     // path delays
     if (A == 1'b1 && B == 1'b1)
       (CI *> S) = (tpllh$CI$S$A_EQ_1_AN_B_EQ_1, tphhl$CI$S$A_EQ_1_AN_B_EQ_1);
     if (A == 1'b1 && B == 1'b0)
       (CI *> S) = (tphlh$CI$S$A_EQ_1_AN_B_EQ_0, tplhl$CI$S$A_EQ_1_AN_B_EQ_0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> S) = (tphlh$CI$S$A_EQ_0_AN_B_EQ_1, tplhl$CI$S$A_EQ_0_AN_B_EQ_1);
     if (A == 1'b0 && B == 1'b0)
       (CI *> S) = (tpllh$CI$S$A_EQ_0_AN_B_EQ_0, tphhl$CI$S$A_EQ_0_AN_B_EQ_0);
     ifnone
       (CI *> S) = (tpllh$CI$S,tplhl$CI$S);

     if (A == 1'b1 && B == 1'b0)
       (CI *> NCO) = (tphlh$CI$NCO$A_EQ_1_AN_B_EQ_0, tplhl$CI$NCO$A_EQ_1_AN_B_EQ_0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> NCO) = (tphlh$CI$NCO$A_EQ_0_AN_B_EQ_1, tplhl$CI$NCO$A_EQ_0_AN_B_EQ_1);
     ifnone
       (CI *> NCO) = (tphlh$CI$NCO,tplhl$CI$NCO);

     if (A == 1'b1 && CI == 1'b1)
       (B *> S) = (tpllh$B$S$A_EQ_1_AN_CI_EQ_1, tphhl$B$S$A_EQ_1_AN_CI_EQ_1);
     if (A == 1'b1 && CI == 1'b0)
       (B *> S) = (tphlh$B$S$A_EQ_1_AN_CI_EQ_0, tplhl$B$S$A_EQ_1_AN_CI_EQ_0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> S) = (tphlh$B$S$A_EQ_0_AN_CI_EQ_1, tplhl$B$S$A_EQ_0_AN_CI_EQ_1);
     if (A == 1'b0 && CI == 1'b0)
       (B *> S) = (tpllh$B$S$A_EQ_0_AN_CI_EQ_0, tphhl$B$S$A_EQ_0_AN_CI_EQ_0);
     ifnone
       (B *> S) = (tpllh$B$S,tplhl$B$S);

     if (A == 1'b1 && CI == 1'b0)
       (B *> NCO) = (tphlh$B$NCO$A_EQ_1_AN_CI_EQ_0, tplhl$B$NCO$A_EQ_1_AN_CI_EQ_0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> NCO) = (tphlh$B$NCO$A_EQ_0_AN_CI_EQ_1, tplhl$B$NCO$A_EQ_0_AN_CI_EQ_1);
     ifnone
       (B *> NCO) = (tphlh$B$NCO,tplhl$B$NCO);

     if (B == 1'b1 && CI == 1'b1)
       (A *> S) = (tpllh$A$S$B_EQ_1_AN_CI_EQ_1, tphhl$A$S$B_EQ_1_AN_CI_EQ_1);
     if (B == 1'b1 && CI == 1'b0)
       (A *> S) = (tphlh$A$S$B_EQ_1_AN_CI_EQ_0, tplhl$A$S$B_EQ_1_AN_CI_EQ_0);
     if (B == 1'b0 && CI == 1'b1)
       (A *> S) = (tphlh$A$S$B_EQ_0_AN_CI_EQ_1, tplhl$A$S$B_EQ_0_AN_CI_EQ_1);
     if (B == 1'b0 && CI == 1'b0)
       (A *> S) = (tpllh$A$S$B_EQ_0_AN_CI_EQ_0, tphhl$A$S$B_EQ_0_AN_CI_EQ_0);
     ifnone
       (A *> S) = (tpllh$A$S,tplhl$A$S);

     if (B == 1'b1 && CI == 1'b0)
       (A *> NCO) = (tphlh$A$NCO$B_EQ_1_AN_CI_EQ_0, tplhl$A$NCO$B_EQ_1_AN_CI_EQ_0);
     if (B == 1'b0 && CI == 1'b1)
       (A *> NCO) = (tphlh$A$NCO$B_EQ_0_AN_CI_EQ_1, tplhl$A$NCO$B_EQ_0_AN_CI_EQ_1);
     ifnone
       (A *> NCO) = (tphlh$A$NCO,tplhl$A$NCO);*/

// path delays
      (posedge A => (NCO +: NCO)) = (1.0, 1.0);
      (negedge A => (NCO -: NCO)) = (1.0, 1.0);
      if (B == 1'b1 && CI == 1'b0) (A -=> NCO) = (1.0, 1.0);
      if (B == 1'b0 && CI == 1'b1) (A -=> NCO) = (1.0, 1.0);
 
      if (B == 1'b1 && CI == 1'b1) (A +=> S) = (1.0, 1.0);
      if (B == 1'b0 && CI == 1'b0) (A +=> S) = (1.0, 1.0);
      if (B == 1'b1 && CI == 1'b0) (A -=> S) = (1.0, 1.0);
      if (B == 1'b0 && CI == 1'b1) (A -=> S) = (1.0, 1.0);

   

      (posedge B => (S +: S)) = (1.0, 1.0);
      (negedge B => (S -: S)) = (1.0, 1.0);
      if (A == 1'b1 && CI == 1'b0) (B -=> NCO) = (1.0, 1.0);
      if (A == 1'b0 && CI == 1'b1) (B -=> NCO) = (1.0, 1.0);
  
      if (A == 1'b1 && CI == 1'b1) (B +=> S) = (1.0, 1.0);
      if (A == 1'b0 && CI == 1'b0) (B +=> S) = (1.0, 1.0);
      if (A == 1'b0 && CI == 1'b1) (B -=> S) = (1.0, 1.0);
      if (A == 1'b1 && CI == 1'b0) (B -=> S) = (1.0, 1.0);
   

      (posedge CI => (S +: S)) = (1.0, 1.0);
      (negedge CI => (S -: S)) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0) (CI +=> NCO) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1) (CI +=> NCO) = (1.0, 1.0);

      if (A == 1'b1 && B == 1'b1) (CI +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b0) (CI +=> S) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0) (CI -=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1) (CI -=> S) = (1.0, 1.0);


   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_FA03D1 (CO, S, A, B, NCI);
input  A ;
input  B ;
input  NCI ;
output CO ;
output S ;

   not (I0_out, NCI);
   and (I1_out, I0_out, A);
   and (I2_out, A, B);
   not (I4_out, NCI);
   and (I5_out, B, I4_out);
   or  (CO, I1_out, I2_out, I5_out);
   xor (I7_out, A, B);
   xor (I8_out, I7_out, NCI);
   not (S, I8_out);

   specify
     // delay parameters
/*     specparam
       tpllh$A$CO = 1.0,
       tphhl$A$CO = 1.0,
       tpllh$A$S = 1.0,
       tplhl$A$S = 1.0,
       tphlh$A$S = 1.0,
       tphhl$A$S = 1.0,
       tpllh$B$CO = 1.0,
       tphhl$B$CO = 1.0,
       tpllh$B$S = 1.0,
       tplhl$B$S = 1.0,
       tphlh$B$S = 1.0,
       tphhl$B$S = 1.0,
       tpllh$NCI$S = 1.0,
       tplhl$NCI$S = 1.0,
       tphlh$NCI$S = 1.0,
       tphhl$NCI$S = 1.0,
       tplhl$NCI$CO = 1.0,
       tphlh$NCI$CO = 1.0,
       tpllh$A$CO$B_EQ_0_AN_NCI_EQ_0 = 1.0,
       tphhl$A$CO$B_EQ_0_AN_NCI_EQ_0 = 1.0,
       tpllh$A$CO$B_EQ_1_AN_NCI_EQ_1 = 1.0,
       tphhl$A$CO$B_EQ_1_AN_NCI_EQ_1 = 1.0,
       tpllh$A$S$B_EQ_1_AN_NCI_EQ_0 = 1.0,
       tphhl$A$S$B_EQ_1_AN_NCI_EQ_0 = 1.0,
       tpllh$A$S$B_EQ_0_AN_NCI_EQ_1 = 1.0,
       tphhl$A$S$B_EQ_0_AN_NCI_EQ_1 = 1.0,
       tplhl$A$S$B_EQ_0_AN_NCI_EQ_0 = 1.0,
       tphlh$A$S$B_EQ_0_AN_NCI_EQ_0 = 1.0,
       tplhl$A$S$B_EQ_1_AN_NCI_EQ_1 = 1.0,
       tphlh$A$S$B_EQ_1_AN_NCI_EQ_1 = 1.0,
       tpllh$B$CO$A_EQ_1_AN_NCI_EQ_1 = 1.0,
       tphhl$B$CO$A_EQ_1_AN_NCI_EQ_1 = 1.0,
       tpllh$B$CO$A_EQ_0_AN_NCI_EQ_0 = 1.0,
       tphhl$B$CO$A_EQ_0_AN_NCI_EQ_0 = 1.0,
       tpllh$B$S$A_EQ_1_AN_NCI_EQ_0 = 1.0,
       tphhl$B$S$A_EQ_1_AN_NCI_EQ_0 = 1.0,
       tpllh$B$S$A_EQ_0_AN_NCI_EQ_1 = 1.0,
       tphhl$B$S$A_EQ_0_AN_NCI_EQ_1 = 1.0,
       tplhl$B$S$A_EQ_1_AN_NCI_EQ_1 = 1.0,
       tphlh$B$S$A_EQ_1_AN_NCI_EQ_1 = 1.0,
       tplhl$B$S$A_EQ_0_AN_NCI_EQ_0 = 1.0,
       tphlh$B$S$A_EQ_0_AN_NCI_EQ_0 = 1.0,
       tpllh$NCI$S$A_EQ_1_AN_B_EQ_0 = 1.0,
       tphhl$NCI$S$A_EQ_1_AN_B_EQ_0 = 1.0,
       tpllh$NCI$S$A_EQ_0_AN_B_EQ_1 = 1.0,
       tphhl$NCI$S$A_EQ_0_AN_B_EQ_1 = 1.0,
       tplhl$NCI$S$A_EQ_1_AN_B_EQ_1 = 1.0,
       tphlh$NCI$S$A_EQ_1_AN_B_EQ_1 = 1.0,
       tplhl$NCI$S$A_EQ_0_AN_B_EQ_0 = 1.0,
       tphlh$NCI$S$A_EQ_0_AN_B_EQ_0 = 1.0,
       tplhl$NCI$CO$A_EQ_1_AN_B_EQ_0 = 1.0,
       tphlh$NCI$CO$A_EQ_1_AN_B_EQ_0 = 1.0,
       tplhl$NCI$CO$A_EQ_0_AN_B_EQ_1 = 1.0,
       tphlh$NCI$CO$A_EQ_0_AN_B_EQ_1 = 1.0;

     // path delays
     if (A == 1'b1 && B == 1'b1)
       (NCI *> S) = (tphlh$NCI$S$A_EQ_1_AN_B_EQ_1, tplhl$NCI$S$A_EQ_1_AN_B_EQ_1);
     if (A == 1'b1 && B == 1'b0)
       (NCI *> S) = (tpllh$NCI$S$A_EQ_1_AN_B_EQ_0, tphhl$NCI$S$A_EQ_1_AN_B_EQ_0);
     if (A == 1'b0 && B == 1'b1)
       (NCI *> S) = (tpllh$NCI$S$A_EQ_0_AN_B_EQ_1, tphhl$NCI$S$A_EQ_0_AN_B_EQ_1);
     if (A == 1'b0 && B == 1'b0)
       (NCI *> S) = (tphlh$NCI$S$A_EQ_0_AN_B_EQ_0, tplhl$NCI$S$A_EQ_0_AN_B_EQ_0);
     ifnone
       (NCI *> S) = (tpllh$NCI$S,tplhl$NCI$S);

     if (A == 1'b1 && B == 1'b0)
       (NCI *> CO) = (tphlh$NCI$CO$A_EQ_1_AN_B_EQ_0, tplhl$NCI$CO$A_EQ_1_AN_B_EQ_0);
     if (A == 1'b0 && B == 1'b1)
       (NCI *> CO) = (tphlh$NCI$CO$A_EQ_0_AN_B_EQ_1, tplhl$NCI$CO$A_EQ_0_AN_B_EQ_1);
     ifnone
       (NCI *> CO) = (tphlh$NCI$CO,tplhl$NCI$CO);

     if (A == 1'b1 && NCI == 1'b1)
       (B *> S) = (tphlh$B$S$A_EQ_1_AN_NCI_EQ_1, tplhl$B$S$A_EQ_1_AN_NCI_EQ_1);
     if (A == 1'b1 && NCI == 1'b0)
       (B *> S) = (tpllh$B$S$A_EQ_1_AN_NCI_EQ_0, tphhl$B$S$A_EQ_1_AN_NCI_EQ_0);
     if (A == 1'b0 && NCI == 1'b1)
       (B *> S) = (tpllh$B$S$A_EQ_0_AN_NCI_EQ_1, tphhl$B$S$A_EQ_0_AN_NCI_EQ_1);
     if (A == 1'b0 && NCI == 1'b0)
       (B *> S) = (tphlh$B$S$A_EQ_0_AN_NCI_EQ_0, tplhl$B$S$A_EQ_0_AN_NCI_EQ_0);
     ifnone
       (B *> S) = (tpllh$B$S,tplhl$B$S);

     if (A == 1'b1 && NCI == 1'b1)
       (B *> CO) = (tpllh$B$CO$A_EQ_1_AN_NCI_EQ_1, tphhl$B$CO$A_EQ_1_AN_NCI_EQ_1);
     if (A == 1'b0 && NCI == 1'b0)
       (B *> CO) = (tpllh$B$CO$A_EQ_0_AN_NCI_EQ_0, tphhl$B$CO$A_EQ_0_AN_NCI_EQ_0);
     ifnone
       (B *> CO) = (tpllh$B$CO,tphhl$B$CO);

     if (B == 1'b1 && NCI == 1'b1)
       (A *> S) = (tphlh$A$S$B_EQ_1_AN_NCI_EQ_1, tplhl$A$S$B_EQ_1_AN_NCI_EQ_1);
     if (B == 1'b1 && NCI == 1'b0)
       (A *> S) = (tpllh$A$S$B_EQ_1_AN_NCI_EQ_0, tphhl$A$S$B_EQ_1_AN_NCI_EQ_0);
     if (B == 1'b0 && NCI == 1'b1)
       (A *> S) = (tpllh$A$S$B_EQ_0_AN_NCI_EQ_1, tphhl$A$S$B_EQ_0_AN_NCI_EQ_1);
     if (B == 1'b0 && NCI == 1'b0)
       (A *> S) = (tphlh$A$S$B_EQ_0_AN_NCI_EQ_0, tplhl$A$S$B_EQ_0_AN_NCI_EQ_0);
     ifnone
       (A *> S) = (tpllh$A$S,tplhl$A$S);

     if (B == 1'b1 && NCI == 1'b1)
       (A *> CO) = (tpllh$A$CO$B_EQ_1_AN_NCI_EQ_1, tphhl$A$CO$B_EQ_1_AN_NCI_EQ_1);
     if (B == 1'b0 && NCI == 1'b0)
       (A *> CO) = (tpllh$A$CO$B_EQ_0_AN_NCI_EQ_0, tphhl$A$CO$B_EQ_0_AN_NCI_EQ_0);
     ifnone
       (A *> CO) = (tpllh$A$CO,tphhl$A$CO);*/

// path delays
      (posedge A => (S +: S)) = (1.0, 1.0);
      (negedge A => (S -: S)) = (1.0, 1.0);
      if (B == 1'b0 && NCI == 1'b0) (A +=> CO) = (1.0, 1.0);
      if (B == 1'b1 && NCI == 1'b1) (A +=> CO) = (1.0, 1.0);
 
      if (B == 1'b1 && NCI == 1'b0) (A +=> S) = (1.0, 1.0);
      if (B == 1'b0 && NCI == 1'b1) (A +=> S) = (1.0, 1.0);
      if (B == 1'b0 && NCI == 1'b0) (A -=> S) = (1.0, 1.0);
      if (B == 1'b1 && NCI == 1'b1) (A -=> S) = (1.0, 1.0);

   

      (posedge B => (S +: S)) = (1.0, 1.0);
      (negedge B => (S -: S)) = (1.0, 1.0);
      if (A == 1'b1 && NCI == 1'b1) (B +=> CO) = (1.0, 1.0);
      if (A == 1'b0 && NCI == 1'b0) (B +=> CO) = (1.0, 1.0);
  
      if (A == 1'b1 && NCI == 1'b0) (B +=> S) = (1.0, 1.0);
      if (A == 1'b0 && NCI == 1'b1) (B +=> S) = (1.0, 1.0);
      if (A == 1'b1 && NCI == 1'b1) (B -=> S) = (1.0, 1.0);
      if (A == 1'b0 && NCI == 1'b0) (B -=> S) = (1.0, 1.0);
   

      (posedge NCI => (S +: S)) = (1.0, 1.0);
      (negedge NCI => (S -: S)) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0) (NCI -=> CO) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1) (NCI -=> CO) = (1.0, 1.0);

      if (A == 1'b1 && B == 1'b0) (NCI +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1) (NCI +=> S) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b1) (NCI -=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b0) (NCI -=> S) = (1.0, 1.0);


   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_FA03D2 (CO, S, A, B, NCI);
input  A ;
input  B ;
input  NCI ;
output CO ;
output S ;

   not (I0_out, NCI);
   and (I1_out, I0_out, A);
   and (I2_out, A, B);
   not (I4_out, NCI);
   and (I5_out, B, I4_out);
   or  (CO, I1_out, I2_out, I5_out);
   xor (I7_out, A, B);
   xor (I8_out, I7_out, NCI);
   not (S, I8_out);

   specify
     // delay parameters
   /*  specparam
       tpllh$A$CO = 1.0,
       tphhl$A$CO = 1.0,
       tpllh$A$S = 1.0,
       tplhl$A$S = 1.0,
       tphlh$A$S = 1.0,
       tphhl$A$S = 1.0,
       tpllh$B$CO = 1.0,
       tphhl$B$CO = 1.0,
       tpllh$B$S = 1.0,
       tplhl$B$S = 1.0,
       tphlh$B$S = 1.0,
       tphhl$B$S = 1.0,
       tpllh$NCI$S = 1.0,
       tplhl$NCI$S = 1.0,
       tphlh$NCI$S = 1.0,
       tphhl$NCI$S = 1.0,
       tplhl$NCI$CO = 1.0,
       tphlh$NCI$CO = 1.0,
       tpllh$A$CO$B_EQ_0_AN_NCI_EQ_0 = 1.0,
       tphhl$A$CO$B_EQ_0_AN_NCI_EQ_0 = 1.0,
       tpllh$A$CO$B_EQ_1_AN_NCI_EQ_1 = 1.0,
       tphhl$A$CO$B_EQ_1_AN_NCI_EQ_1 = 1.0,
       tpllh$A$S$B_EQ_1_AN_NCI_EQ_0 = 1.0,
       tphhl$A$S$B_EQ_1_AN_NCI_EQ_0 = 1.0,
       tpllh$A$S$B_EQ_0_AN_NCI_EQ_1 = 1.0,
       tphhl$A$S$B_EQ_0_AN_NCI_EQ_1 = 1.0,
       tplhl$A$S$B_EQ_0_AN_NCI_EQ_0 = 1.0,
       tphlh$A$S$B_EQ_0_AN_NCI_EQ_0 = 1.0,
       tplhl$A$S$B_EQ_1_AN_NCI_EQ_1 = 1.0,
       tphlh$A$S$B_EQ_1_AN_NCI_EQ_1 = 1.0,
       tpllh$B$CO$A_EQ_1_AN_NCI_EQ_1 = 1.0,
       tphhl$B$CO$A_EQ_1_AN_NCI_EQ_1 = 1.0,
       tpllh$B$CO$A_EQ_0_AN_NCI_EQ_0 = 1.0,
       tphhl$B$CO$A_EQ_0_AN_NCI_EQ_0 = 1.0,
       tpllh$B$S$A_EQ_1_AN_NCI_EQ_0 = 1.0,
       tphhl$B$S$A_EQ_1_AN_NCI_EQ_0 = 1.0,
       tpllh$B$S$A_EQ_0_AN_NCI_EQ_1 = 1.0,
       tphhl$B$S$A_EQ_0_AN_NCI_EQ_1 = 1.0,
       tplhl$B$S$A_EQ_1_AN_NCI_EQ_1 = 1.0,
       tphlh$B$S$A_EQ_1_AN_NCI_EQ_1 = 1.0,
       tplhl$B$S$A_EQ_0_AN_NCI_EQ_0 = 1.0,
       tphlh$B$S$A_EQ_0_AN_NCI_EQ_0 = 1.0,
       tpllh$NCI$S$A_EQ_1_AN_B_EQ_0 = 1.0,
       tphhl$NCI$S$A_EQ_1_AN_B_EQ_0 = 1.0,
       tpllh$NCI$S$A_EQ_0_AN_B_EQ_1 = 1.0,
       tphhl$NCI$S$A_EQ_0_AN_B_EQ_1 = 1.0,
       tplhl$NCI$S$A_EQ_1_AN_B_EQ_1 = 1.0,
       tphlh$NCI$S$A_EQ_1_AN_B_EQ_1 = 1.0,
       tplhl$NCI$S$A_EQ_0_AN_B_EQ_0 = 1.0,
       tphlh$NCI$S$A_EQ_0_AN_B_EQ_0 = 1.0,
       tplhl$NCI$CO$A_EQ_1_AN_B_EQ_0 = 1.0,
       tphlh$NCI$CO$A_EQ_1_AN_B_EQ_0 = 1.0,
       tplhl$NCI$CO$A_EQ_0_AN_B_EQ_1 = 1.0,
       tphlh$NCI$CO$A_EQ_0_AN_B_EQ_1 = 1.0;

     // path delays
     if (A == 1'b1 && B == 1'b1)
       (NCI *> S) = (tphlh$NCI$S$A_EQ_1_AN_B_EQ_1, tplhl$NCI$S$A_EQ_1_AN_B_EQ_1);
     if (A == 1'b1 && B == 1'b0)
       (NCI *> S) = (tpllh$NCI$S$A_EQ_1_AN_B_EQ_0, tphhl$NCI$S$A_EQ_1_AN_B_EQ_0);
     if (A == 1'b0 && B == 1'b1)
       (NCI *> S) = (tpllh$NCI$S$A_EQ_0_AN_B_EQ_1, tphhl$NCI$S$A_EQ_0_AN_B_EQ_1);
     if (A == 1'b0 && B == 1'b0)
       (NCI *> S) = (tphlh$NCI$S$A_EQ_0_AN_B_EQ_0, tplhl$NCI$S$A_EQ_0_AN_B_EQ_0);
     ifnone
       (NCI *> S) = (tpllh$NCI$S,tplhl$NCI$S);

     if (A == 1'b1 && B == 1'b0)
       (NCI *> CO) = (tphlh$NCI$CO$A_EQ_1_AN_B_EQ_0, tplhl$NCI$CO$A_EQ_1_AN_B_EQ_0);
     if (A == 1'b0 && B == 1'b1)
       (NCI *> CO) = (tphlh$NCI$CO$A_EQ_0_AN_B_EQ_1, tplhl$NCI$CO$A_EQ_0_AN_B_EQ_1);
     ifnone
       (NCI *> CO) = (tphlh$NCI$CO,tplhl$NCI$CO);

     if (A == 1'b1 && NCI == 1'b1)
       (B *> S) = (tphlh$B$S$A_EQ_1_AN_NCI_EQ_1, tplhl$B$S$A_EQ_1_AN_NCI_EQ_1);
     if (A == 1'b1 && NCI == 1'b0)
       (B *> S) = (tpllh$B$S$A_EQ_1_AN_NCI_EQ_0, tphhl$B$S$A_EQ_1_AN_NCI_EQ_0);
     if (A == 1'b0 && NCI == 1'b1)
       (B *> S) = (tpllh$B$S$A_EQ_0_AN_NCI_EQ_1, tphhl$B$S$A_EQ_0_AN_NCI_EQ_1);
     if (A == 1'b0 && NCI == 1'b0)
       (B *> S) = (tphlh$B$S$A_EQ_0_AN_NCI_EQ_0, tplhl$B$S$A_EQ_0_AN_NCI_EQ_0);
     ifnone
       (B *> S) = (tpllh$B$S,tplhl$B$S);

     if (A == 1'b1 && NCI == 1'b1)
       (B *> CO) = (tpllh$B$CO$A_EQ_1_AN_NCI_EQ_1, tphhl$B$CO$A_EQ_1_AN_NCI_EQ_1);
     if (A == 1'b0 && NCI == 1'b0)
       (B *> CO) = (tpllh$B$CO$A_EQ_0_AN_NCI_EQ_0, tphhl$B$CO$A_EQ_0_AN_NCI_EQ_0);
     ifnone
       (B *> CO) = (tpllh$B$CO,tphhl$B$CO);

     if (B == 1'b1 && NCI == 1'b1)
       (A *> S) = (tphlh$A$S$B_EQ_1_AN_NCI_EQ_1, tplhl$A$S$B_EQ_1_AN_NCI_EQ_1);
     if (B == 1'b1 && NCI == 1'b0)
       (A *> S) = (tpllh$A$S$B_EQ_1_AN_NCI_EQ_0, tphhl$A$S$B_EQ_1_AN_NCI_EQ_0);
     if (B == 1'b0 && NCI == 1'b1)
       (A *> S) = (tpllh$A$S$B_EQ_0_AN_NCI_EQ_1, tphhl$A$S$B_EQ_0_AN_NCI_EQ_1);
     if (B == 1'b0 && NCI == 1'b0)
       (A *> S) = (tphlh$A$S$B_EQ_0_AN_NCI_EQ_0, tplhl$A$S$B_EQ_0_AN_NCI_EQ_0);
     ifnone
       (A *> S) = (tpllh$A$S,tplhl$A$S);

     if (B == 1'b1 && NCI == 1'b1)
       (A *> CO) = (tpllh$A$CO$B_EQ_1_AN_NCI_EQ_1, tphhl$A$CO$B_EQ_1_AN_NCI_EQ_1);
     if (B == 1'b0 && NCI == 1'b0)
       (A *> CO) = (tpllh$A$CO$B_EQ_0_AN_NCI_EQ_0, tphhl$A$CO$B_EQ_0_AN_NCI_EQ_0);
     ifnone
       (A *> CO) = (tpllh$A$CO,tphhl$A$CO);*/

// path delays
      (posedge A => (S +: S)) = (1.0, 1.0);
      (negedge A => (S -: S)) = (1.0, 1.0);
      if (B == 1'b0 && NCI == 1'b0) (A +=> CO) = (1.0, 1.0);
      if (B == 1'b1 && NCI == 1'b1) (A +=> CO) = (1.0, 1.0);
 
      if (B == 1'b1 && NCI == 1'b0) (A +=> S) = (1.0, 1.0);
      if (B == 1'b0 && NCI == 1'b1) (A +=> S) = (1.0, 1.0);
      if (B == 1'b0 && NCI == 1'b0) (A -=> S) = (1.0, 1.0);
      if (B == 1'b1 && NCI == 1'b1) (A -=> S) = (1.0, 1.0);

   

      (posedge B => (S +: S)) = (1.0, 1.0);
      (negedge B => (S -: S)) = (1.0, 1.0);
      if (A == 1'b1 && NCI == 1'b1) (B +=> CO) = (1.0, 1.0);
      if (A == 1'b0 && NCI == 1'b0) (B +=> CO) = (1.0, 1.0);
  
      if (A == 1'b1 && NCI == 1'b0) (B +=> S) = (1.0, 1.0);
      if (A == 1'b0 && NCI == 1'b1) (B +=> S) = (1.0, 1.0);
      if (A == 1'b1 && NCI == 1'b1) (B -=> S) = (1.0, 1.0);
      if (A == 1'b0 && NCI == 1'b0) (B -=> S) = (1.0, 1.0);
   

      (posedge NCI => (S +: S)) = (1.0, 1.0);
      (negedge NCI => (S -: S)) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0) (NCI -=> CO) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1) (NCI -=> CO) = (1.0, 1.0);

      if (A == 1'b1 && B == 1'b0) (NCI +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1) (NCI +=> S) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b1) (NCI -=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b0) (NCI -=> S) = (1.0, 1.0);



   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_FA03D4 (CO, S, A, B, NCI);
input  A ;
input  B ;
input  NCI ;
output CO ;
output S ;

   not (I0_out, NCI);
   and (I1_out, I0_out, A);
   and (I2_out, A, B);
   not (I4_out, NCI);
   and (I5_out, B, I4_out);
   or  (CO, I1_out, I2_out, I5_out);
   xor (I7_out, A, B);
   xor (I8_out, I7_out, NCI);
   not (S, I8_out);

   specify
     // delay parameters
  /*   specparam
       tpllh$A$CO = 1.0,
       tphhl$A$CO = 1.0,
       tpllh$A$S = 1.0,
       tplhl$A$S = 1.0,
       tphlh$A$S = 1.0,
       tphhl$A$S = 1.0,
       tpllh$B$CO = 1.0,
       tphhl$B$CO = 1.0,
       tpllh$B$S = 1.0,
       tplhl$B$S = 1.0,
       tphlh$B$S = 1.0,
       tphhl$B$S = 1.0,
       tpllh$NCI$S = 1.0,
       tplhl$NCI$S = 1.0,
       tphlh$NCI$S = 1.0,
       tphhl$NCI$S = 1.0,
       tplhl$NCI$CO = 1.0,
       tphlh$NCI$CO = 1.0,
       tpllh$A$CO$B_EQ_0_AN_NCI_EQ_0 = 1.0,
       tphhl$A$CO$B_EQ_0_AN_NCI_EQ_0 = 1.0,
       tpllh$A$CO$B_EQ_1_AN_NCI_EQ_1 = 1.0,
       tphhl$A$CO$B_EQ_1_AN_NCI_EQ_1 = 1.0,
       tpllh$A$S$B_EQ_1_AN_NCI_EQ_0 = 1.0,
       tphhl$A$S$B_EQ_1_AN_NCI_EQ_0 = 1.0,
       tpllh$A$S$B_EQ_0_AN_NCI_EQ_1 = 1.0,
       tphhl$A$S$B_EQ_0_AN_NCI_EQ_1 = 1.0,
       tplhl$A$S$B_EQ_0_AN_NCI_EQ_0 = 1.0,
       tphlh$A$S$B_EQ_0_AN_NCI_EQ_0 = 1.0,
       tplhl$A$S$B_EQ_1_AN_NCI_EQ_1 = 1.0,
       tphlh$A$S$B_EQ_1_AN_NCI_EQ_1 = 1.0,
       tpllh$B$CO$A_EQ_1_AN_NCI_EQ_1 = 1.0,
       tphhl$B$CO$A_EQ_1_AN_NCI_EQ_1 = 1.0,
       tpllh$B$CO$A_EQ_0_AN_NCI_EQ_0 = 1.0,
       tphhl$B$CO$A_EQ_0_AN_NCI_EQ_0 = 1.0,
       tpllh$B$S$A_EQ_1_AN_NCI_EQ_0 = 1.0,
       tphhl$B$S$A_EQ_1_AN_NCI_EQ_0 = 1.0,
       tpllh$B$S$A_EQ_0_AN_NCI_EQ_1 = 1.0,
       tphhl$B$S$A_EQ_0_AN_NCI_EQ_1 = 1.0,
       tplhl$B$S$A_EQ_1_AN_NCI_EQ_1 = 1.0,
       tphlh$B$S$A_EQ_1_AN_NCI_EQ_1 = 1.0,
       tplhl$B$S$A_EQ_0_AN_NCI_EQ_0 = 1.0,
       tphlh$B$S$A_EQ_0_AN_NCI_EQ_0 = 1.0,
       tpllh$NCI$S$A_EQ_1_AN_B_EQ_0 = 1.0,
       tphhl$NCI$S$A_EQ_1_AN_B_EQ_0 = 1.0,
       tpllh$NCI$S$A_EQ_0_AN_B_EQ_1 = 1.0,
       tphhl$NCI$S$A_EQ_0_AN_B_EQ_1 = 1.0,
       tplhl$NCI$S$A_EQ_1_AN_B_EQ_1 = 1.0,
       tphlh$NCI$S$A_EQ_1_AN_B_EQ_1 = 1.0,
       tplhl$NCI$S$A_EQ_0_AN_B_EQ_0 = 1.0,
       tphlh$NCI$S$A_EQ_0_AN_B_EQ_0 = 1.0,
       tplhl$NCI$CO$A_EQ_1_AN_B_EQ_0 = 1.0,
       tphlh$NCI$CO$A_EQ_1_AN_B_EQ_0 = 1.0,
       tplhl$NCI$CO$A_EQ_0_AN_B_EQ_1 = 1.0,
       tphlh$NCI$CO$A_EQ_0_AN_B_EQ_1 = 1.0;

     // path delays
     if (A == 1'b1 && B == 1'b1)
       (NCI *> S) = (tphlh$NCI$S$A_EQ_1_AN_B_EQ_1, tplhl$NCI$S$A_EQ_1_AN_B_EQ_1);
     if (A == 1'b1 && B == 1'b0)
       (NCI *> S) = (tpllh$NCI$S$A_EQ_1_AN_B_EQ_0, tphhl$NCI$S$A_EQ_1_AN_B_EQ_0);
     if (A == 1'b0 && B == 1'b1)
       (NCI *> S) = (tpllh$NCI$S$A_EQ_0_AN_B_EQ_1, tphhl$NCI$S$A_EQ_0_AN_B_EQ_1);
     if (A == 1'b0 && B == 1'b0)
       (NCI *> S) = (tphlh$NCI$S$A_EQ_0_AN_B_EQ_0, tplhl$NCI$S$A_EQ_0_AN_B_EQ_0);
     ifnone
       (NCI *> S) = (tpllh$NCI$S,tplhl$NCI$S);

     if (A == 1'b1 && B == 1'b0)
       (NCI *> CO) = (tphlh$NCI$CO$A_EQ_1_AN_B_EQ_0, tplhl$NCI$CO$A_EQ_1_AN_B_EQ_0);
     if (A == 1'b0 && B == 1'b1)
       (NCI *> CO) = (tphlh$NCI$CO$A_EQ_0_AN_B_EQ_1, tplhl$NCI$CO$A_EQ_0_AN_B_EQ_1);
     ifnone
       (NCI *> CO) = (tphlh$NCI$CO,tplhl$NCI$CO);

     if (A == 1'b1 && NCI == 1'b1)
       (B *> S) = (tphlh$B$S$A_EQ_1_AN_NCI_EQ_1, tplhl$B$S$A_EQ_1_AN_NCI_EQ_1);
     if (A == 1'b1 && NCI == 1'b0)
       (B *> S) = (tpllh$B$S$A_EQ_1_AN_NCI_EQ_0, tphhl$B$S$A_EQ_1_AN_NCI_EQ_0);
     if (A == 1'b0 && NCI == 1'b1)
       (B *> S) = (tpllh$B$S$A_EQ_0_AN_NCI_EQ_1, tphhl$B$S$A_EQ_0_AN_NCI_EQ_1);
     if (A == 1'b0 && NCI == 1'b0)
       (B *> S) = (tphlh$B$S$A_EQ_0_AN_NCI_EQ_0, tplhl$B$S$A_EQ_0_AN_NCI_EQ_0);
     ifnone
       (B *> S) = (tpllh$B$S,tplhl$B$S);

     if (A == 1'b1 && NCI == 1'b1)
       (B *> CO) = (tpllh$B$CO$A_EQ_1_AN_NCI_EQ_1, tphhl$B$CO$A_EQ_1_AN_NCI_EQ_1);
     if (A == 1'b0 && NCI == 1'b0)
       (B *> CO) = (tpllh$B$CO$A_EQ_0_AN_NCI_EQ_0, tphhl$B$CO$A_EQ_0_AN_NCI_EQ_0);
     ifnone
       (B *> CO) = (tpllh$B$CO,tphhl$B$CO);

     if (B == 1'b1 && NCI == 1'b1)
       (A *> S) = (tphlh$A$S$B_EQ_1_AN_NCI_EQ_1, tplhl$A$S$B_EQ_1_AN_NCI_EQ_1);
     if (B == 1'b1 && NCI == 1'b0)
       (A *> S) = (tpllh$A$S$B_EQ_1_AN_NCI_EQ_0, tphhl$A$S$B_EQ_1_AN_NCI_EQ_0);
     if (B == 1'b0 && NCI == 1'b1)
       (A *> S) = (tpllh$A$S$B_EQ_0_AN_NCI_EQ_1, tphhl$A$S$B_EQ_0_AN_NCI_EQ_1);
     if (B == 1'b0 && NCI == 1'b0)
       (A *> S) = (tphlh$A$S$B_EQ_0_AN_NCI_EQ_0, tplhl$A$S$B_EQ_0_AN_NCI_EQ_0);
     ifnone
       (A *> S) = (tpllh$A$S,tplhl$A$S);

     if (B == 1'b1 && NCI == 1'b1)
       (A *> CO) = (tpllh$A$CO$B_EQ_1_AN_NCI_EQ_1, tphhl$A$CO$B_EQ_1_AN_NCI_EQ_1);
     if (B == 1'b0 && NCI == 1'b0)
       (A *> CO) = (tpllh$A$CO$B_EQ_0_AN_NCI_EQ_0, tphhl$A$CO$B_EQ_0_AN_NCI_EQ_0);
     ifnone
       (A *> CO) = (tpllh$A$CO,tphhl$A$CO);*/

// path delays
      (posedge A => (CO +: CO)) = (1.0, 1.0);
      (negedge A => (CO -: CO)) = (1.0, 1.0);
      if (B == 1'b0 && NCI == 1'b0) (A +=> CO) = (1.0, 1.0);
      if (B == 1'b1 && NCI == 1'b1) (A +=> CO) = (1.0, 1.0);
 
      if (B == 1'b1 && NCI == 1'b0) (A +=> S) = (1.0, 1.0);
      if (B == 1'b0 && NCI == 1'b1) (A +=> S) = (1.0, 1.0);
      if (B == 1'b0 && NCI == 1'b0) (A -=> S) = (1.0, 1.0);
      if (B == 1'b1 && NCI == 1'b1) (A -=> S) = (1.0, 1.0);

   

      (posedge B => (S +: S)) = (1.0, 1.0);
      (negedge B => (S -: S)) = (1.0, 1.0);
      if (A == 1'b1 && NCI == 1'b1) (B +=> CO) = (1.0, 1.0);
      if (A == 1'b0 && NCI == 1'b0) (B +=> CO) = (1.0, 1.0);
  
      if (A == 1'b1 && NCI == 1'b0) (B +=> S) = (1.0, 1.0);
      if (A == 1'b0 && NCI == 1'b1) (B +=> S) = (1.0, 1.0);
      if (A == 1'b1 && NCI == 1'b1) (B -=> S) = (1.0, 1.0);
      if (A == 1'b0 && NCI == 1'b0) (B -=> S) = (1.0, 1.0);
   

      (posedge NCI => (S +: S)) = (1.0, 1.0);
      (negedge NCI => (S -: S)) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0) (NCI -=> CO) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1) (NCI -=> CO) = (1.0, 1.0);

      if (A == 1'b1 && B == 1'b0) (NCI +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1) (NCI +=> S) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b1) (NCI -=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b0) (NCI -=> S) = (1.0, 1.0);



   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_FA04D1 (NCO1, NCO2, S, A, B, CI1, CI2, CS);
input  A ;
input  B ;
input  CI1 ;
input  CI2 ;
input  CS ;
output NCO1 ;
output NCO2 ;
output S ;

   and (I0_out, A, B);
   and (I1_out, B, CI1);
   and (I3_out, CI1, A);
   or  (I4_out, I0_out, I1_out, I3_out);
   not (NCO1, I4_out);
   and (I6_out, A, B);
   and (I7_out, B, CI2);
   and (I9_out, CI2, A);
   or  (I10_out, I6_out, I7_out, I9_out);
   not (NCO2, I10_out);
   udp_mux2 (I12_out, CI1, CI2, CS);
   xor (I13_out, I12_out, A);
   xor (S, I13_out, B);

   specify
     // delay parameters
   /*  specparam
       tpllh$A$S = 1.0,
       tplhl$A$S = 1.0,
       tphlh$A$S = 1.0,
       tphhl$A$S = 1.0,
       tplhl$A$NCO2 = 1.0,
       tphlh$A$NCO2 = 1.0,
       tplhl$A$NCO1 = 1.0,
       tphlh$A$NCO1 = 1.0,
       tpllh$B$S = 1.0,
       tplhl$B$S = 1.0,
       tphlh$B$S = 1.0,
       tphhl$B$S = 1.0,
       tplhl$B$NCO2 = 1.0,
       tphlh$B$NCO2 = 1.0,
       tplhl$B$NCO1 = 1.0,
       tphlh$B$NCO1 = 1.0,
       tpllh$CI1$S = 1.0,
       tplhl$CI1$S = 1.0,
       tphlh$CI1$S = 1.0,
       tphhl$CI1$S = 1.0,
       tplhl$CI1$NCO1 = 1.0,
       tphlh$CI1$NCO1 = 1.0,
       tpllh$CI2$S = 1.0,
       tplhl$CI2$S = 1.0,
       tphlh$CI2$S = 1.0,
       tphhl$CI2$S = 1.0,
       tplhl$CI2$NCO2 = 1.0,
       tphlh$CI2$NCO2 = 1.0,
       tpllh$CS$S = 1.0,
       tplhl$CS$S = 1.0,
       tphlh$CS$S = 1.0,
       tphhl$CS$S = 1.0,
       tpllh$A$S$B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tphhl$A$S$B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tpllh$A$S$B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tphhl$A$S$B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tpllh$A$S$B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tphhl$A$S$B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tpllh$A$S$B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tphhl$A$S$B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tpllh$A$S$B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1 = 1.0,
       tphhl$A$S$B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1 = 1.0,
       tpllh$A$S$B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tphhl$A$S$B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tplhl$A$S$B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tphlh$A$S$B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tplhl$A$S$B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tphlh$A$S$B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tplhl$A$S$B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1 = 1.0,
       tphlh$A$S$B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1 = 1.0,
       tplhl$A$S$B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tphlh$A$S$B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tplhl$A$S$B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tphlh$A$S$B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tplhl$A$S$B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tphlh$A$S$B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tplhl$A$NCO2$B_EQ_1_AN_CI2_EQ_0 = 1.0,
       tphlh$A$NCO2$B_EQ_1_AN_CI2_EQ_0 = 1.0,
       tplhl$A$NCO2$B_EQ_0_AN_CI2_EQ_1 = 1.0,
       tphlh$A$NCO2$B_EQ_0_AN_CI2_EQ_1 = 1.0,
       tplhl$A$NCO1$B_EQ_1_AN_CI1_EQ_0 = 1.0,
       tphlh$A$NCO1$B_EQ_1_AN_CI1_EQ_0 = 1.0,
       tplhl$A$NCO1$B_EQ_0_AN_CI1_EQ_1 = 1.0,
       tphlh$A$NCO1$B_EQ_0_AN_CI1_EQ_1 = 1.0,
       tpllh$B$S$A_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tphhl$B$S$A_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tpllh$B$S$A_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tphhl$B$S$A_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tpllh$B$S$A_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tphhl$B$S$A_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tpllh$B$S$A_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1 = 1.0,
       tphhl$B$S$A_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1 = 1.0,
       tpllh$B$S$A_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tphhl$B$S$A_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tpllh$B$S$A_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tphhl$B$S$A_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tplhl$B$S$A_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tphlh$B$S$A_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tplhl$B$S$A_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tphlh$B$S$A_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tplhl$B$S$A_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1 = 1.0,
       tphlh$B$S$A_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1 = 1.0,
       tplhl$B$S$A_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tphlh$B$S$A_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tplhl$B$S$A_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tphlh$B$S$A_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tplhl$B$S$A_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tphlh$B$S$A_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tplhl$B$NCO2$A_EQ_1_AN_CI2_EQ_0 = 1.0,
       tphlh$B$NCO2$A_EQ_1_AN_CI2_EQ_0 = 1.0,
       tplhl$B$NCO2$A_EQ_0_AN_CI2_EQ_1 = 1.0,
       tphlh$B$NCO2$A_EQ_0_AN_CI2_EQ_1 = 1.0,
       tplhl$B$NCO1$A_EQ_1_AN_CI1_EQ_0 = 1.0,
       tphlh$B$NCO1$A_EQ_1_AN_CI1_EQ_0 = 1.0,
       tplhl$B$NCO1$A_EQ_0_AN_CI1_EQ_1 = 1.0,
       tphlh$B$NCO1$A_EQ_0_AN_CI1_EQ_1 = 1.0,
       tpllh$CI1$S$A_EQ_1_AN_B_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tphhl$CI1$S$A_EQ_1_AN_B_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tpllh$CI1$S$A_EQ_0_AN_B_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tphhl$CI1$S$A_EQ_0_AN_B_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tplhl$CI1$S$A_EQ_1_AN_B_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tphlh$CI1$S$A_EQ_1_AN_B_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tplhl$CI1$S$A_EQ_0_AN_B_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tphlh$CI1$S$A_EQ_0_AN_B_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tplhl$CI1$S$A_EQ_1_AN_B_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tphlh$CI1$S$A_EQ_1_AN_B_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tplhl$CI1$S$A_EQ_0_AN_B_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tphlh$CI1$S$A_EQ_0_AN_B_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tplhl$CI1$NCO1$A_EQ_0_AN_B_EQ_1 = 1.0,
       tphlh$CI1$NCO1$A_EQ_0_AN_B_EQ_1 = 1.0,
       tplhl$CI1$NCO1$A_EQ_1_AN_B_EQ_0 = 1.0,
       tphlh$CI1$NCO1$A_EQ_1_AN_B_EQ_0 = 1.0,
       tpllh$CI2$S$A_EQ_1_AN_B_EQ_1_AN_CI1_EQ_1_AN_CS_EQ_1 = 1.0,
       tphhl$CI2$S$A_EQ_1_AN_B_EQ_1_AN_CI1_EQ_1_AN_CS_EQ_1 = 1.0,
       tpllh$CI2$S$A_EQ_0_AN_B_EQ_0_AN_CI1_EQ_0_AN_CS_EQ_1 = 1.0,
       tphhl$CI2$S$A_EQ_0_AN_B_EQ_0_AN_CI1_EQ_0_AN_CS_EQ_1 = 1.0,
       tplhl$CI2$S$A_EQ_0_AN_B_EQ_1_AN_CI1_EQ_0_AN_CS_EQ_1 = 1.0,
       tphlh$CI2$S$A_EQ_0_AN_B_EQ_1_AN_CI1_EQ_0_AN_CS_EQ_1 = 1.0,
       tplhl$CI2$S$A_EQ_1_AN_B_EQ_0_AN_CI1_EQ_0_AN_CS_EQ_1 = 1.0,
       tphlh$CI2$S$A_EQ_1_AN_B_EQ_0_AN_CI1_EQ_0_AN_CS_EQ_1 = 1.0,
       tplhl$CI2$S$A_EQ_0_AN_B_EQ_1_AN_CI1_EQ_1_AN_CS_EQ_1 = 1.0,
       tphlh$CI2$S$A_EQ_0_AN_B_EQ_1_AN_CI1_EQ_1_AN_CS_EQ_1 = 1.0,
       tplhl$CI2$S$A_EQ_1_AN_B_EQ_0_AN_CI1_EQ_1_AN_CS_EQ_1 = 1.0,
       tphlh$CI2$S$A_EQ_1_AN_B_EQ_0_AN_CI1_EQ_1_AN_CS_EQ_1 = 1.0,
       tplhl$CI2$NCO2$A_EQ_0_AN_B_EQ_1 = 1.0,
       tphlh$CI2$NCO2$A_EQ_0_AN_B_EQ_1 = 1.0,
       tplhl$CI2$NCO2$A_EQ_1_AN_B_EQ_0 = 1.0,
       tphlh$CI2$NCO2$A_EQ_1_AN_B_EQ_0 = 1.0,
       tpllh$CS$S$A_EQ_1_AN_B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1 = 1.0,
       tphhl$CS$S$A_EQ_1_AN_B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1 = 1.0,
       tpllh$CS$S$A_EQ_0_AN_B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1 = 1.0,
       tphhl$CS$S$A_EQ_0_AN_B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1 = 1.0,
       tplhl$CS$S$A_EQ_1_AN_B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0 = 1.0,
       tphlh$CS$S$A_EQ_1_AN_B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0 = 1.0,
       tplhl$CS$S$A_EQ_0_AN_B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0 = 1.0,
       tphlh$CS$S$A_EQ_0_AN_B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0 = 1.0;

     // path delays
     if (A == 1'b1 && B == 1'b1 && CI1 == 1'b1 && CI2 == 1'b0)
       (CS *> S) = (tphlh$CS$S$A_EQ_1_AN_B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0, tplhl$CS$S$A_EQ_1_AN_B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0);
     if (A == 1'b1 && B == 1'b1 && CI1 == 1'b0 && CI2 == 1'b1)
       (CS *> S) = (tpllh$CS$S$A_EQ_1_AN_B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1, tphhl$CS$S$A_EQ_1_AN_B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1);
     if (A == 1'b0 && B == 1'b0 && CI1 == 1'b1 && CI2 == 1'b0)
       (CS *> S) = (tphlh$CS$S$A_EQ_0_AN_B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0, tplhl$CS$S$A_EQ_0_AN_B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0);
     if (A == 1'b0 && B == 1'b0 && CI1 == 1'b0 && CI2 == 1'b1)
       (CS *> S) = (tpllh$CS$S$A_EQ_0_AN_B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1, tphhl$CS$S$A_EQ_0_AN_B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1);
     ifnone
       (CS *> S) = (tpllh$CS$S,tplhl$CS$S);

     if (A == 1'b1 && B == 1'b1 && CI1 == 1'b1 && CS == 1'b1)
       (CI2 *> S) = (tpllh$CI2$S$A_EQ_1_AN_B_EQ_1_AN_CI1_EQ_1_AN_CS_EQ_1, tphhl$CI2$S$A_EQ_1_AN_B_EQ_1_AN_CI1_EQ_1_AN_CS_EQ_1);
     if (A == 1'b1 && B == 1'b0 && CI1 == 1'b1 && CS == 1'b1)
       (CI2 *> S) = (tphlh$CI2$S$A_EQ_1_AN_B_EQ_0_AN_CI1_EQ_1_AN_CS_EQ_1, tplhl$CI2$S$A_EQ_1_AN_B_EQ_0_AN_CI1_EQ_1_AN_CS_EQ_1);
     if (A == 1'b1 && B == 1'b0 && CI1 == 1'b0 && CS == 1'b1)
       (CI2 *> S) = (tphlh$CI2$S$A_EQ_1_AN_B_EQ_0_AN_CI1_EQ_0_AN_CS_EQ_1, tplhl$CI2$S$A_EQ_1_AN_B_EQ_0_AN_CI1_EQ_0_AN_CS_EQ_1);
     if (A == 1'b0 && B == 1'b1 && CI1 == 1'b1 && CS == 1'b1)
       (CI2 *> S) = (tphlh$CI2$S$A_EQ_0_AN_B_EQ_1_AN_CI1_EQ_1_AN_CS_EQ_1, tplhl$CI2$S$A_EQ_0_AN_B_EQ_1_AN_CI1_EQ_1_AN_CS_EQ_1);
     if (A == 1'b0 && B == 1'b1 && CI1 == 1'b0 && CS == 1'b1)
       (CI2 *> S) = (tphlh$CI2$S$A_EQ_0_AN_B_EQ_1_AN_CI1_EQ_0_AN_CS_EQ_1, tplhl$CI2$S$A_EQ_0_AN_B_EQ_1_AN_CI1_EQ_0_AN_CS_EQ_1);
     if (A == 1'b0 && B == 1'b0 && CI1 == 1'b0 && CS == 1'b1)
       (CI2 *> S) = (tpllh$CI2$S$A_EQ_0_AN_B_EQ_0_AN_CI1_EQ_0_AN_CS_EQ_1, tphhl$CI2$S$A_EQ_0_AN_B_EQ_0_AN_CI1_EQ_0_AN_CS_EQ_1);
     ifnone
       (CI2 *> S) = (tpllh$CI2$S,tplhl$CI2$S);

     if (A == 1'b1 && B == 1'b0)
       (CI2 *> NCO2) = (tphlh$CI2$NCO2$A_EQ_1_AN_B_EQ_0, tplhl$CI2$NCO2$A_EQ_1_AN_B_EQ_0);
     if (A == 1'b0 && B == 1'b1)
       (CI2 *> NCO2) = (tphlh$CI2$NCO2$A_EQ_0_AN_B_EQ_1, tplhl$CI2$NCO2$A_EQ_0_AN_B_EQ_1);
     ifnone
       (CI2 *> NCO2) = (tphlh$CI2$NCO2,tplhl$CI2$NCO2);

     if (A == 1'b1 && B == 1'b1 && CI2 == 1'b1 && CS == 1'b0)
       (CI1 *> S) = (tpllh$CI1$S$A_EQ_1_AN_B_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_0, tphhl$CI1$S$A_EQ_1_AN_B_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_0);
     if (A == 1'b1 && B == 1'b0 && CI2 == 1'b1 && CS == 1'b0)
       (CI1 *> S) = (tphlh$CI1$S$A_EQ_1_AN_B_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0, tplhl$CI1$S$A_EQ_1_AN_B_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0);
     if (A == 1'b1 && B == 1'b0 && CI2 == 1'b0 && CS == 1'b0)
       (CI1 *> S) = (tphlh$CI1$S$A_EQ_1_AN_B_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0, tplhl$CI1$S$A_EQ_1_AN_B_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0);
     if (A == 1'b0 && B == 1'b1 && CI2 == 1'b1 && CS == 1'b0)
       (CI1 *> S) = (tphlh$CI1$S$A_EQ_0_AN_B_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_0, tplhl$CI1$S$A_EQ_0_AN_B_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_0);
     if (A == 1'b0 && B == 1'b1 && CI2 == 1'b0 && CS == 1'b0)
       (CI1 *> S) = (tphlh$CI1$S$A_EQ_0_AN_B_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0, tplhl$CI1$S$A_EQ_0_AN_B_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0);
     if (A == 1'b0 && B == 1'b0 && CI2 == 1'b0 && CS == 1'b0)
       (CI1 *> S) = (tpllh$CI1$S$A_EQ_0_AN_B_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0, tphhl$CI1$S$A_EQ_0_AN_B_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0);
     ifnone
       (CI1 *> S) = (tpllh$CI1$S,tplhl$CI1$S);

     if (A == 1'b1 && B == 1'b0)
       (CI1 *> NCO1) = (tphlh$CI1$NCO1$A_EQ_1_AN_B_EQ_0, tplhl$CI1$NCO1$A_EQ_1_AN_B_EQ_0);
     if (A == 1'b0 && B == 1'b1)
       (CI1 *> NCO1) = (tphlh$CI1$NCO1$A_EQ_0_AN_B_EQ_1, tplhl$CI1$NCO1$A_EQ_0_AN_B_EQ_1);
     ifnone
       (CI1 *> NCO1) = (tphlh$CI1$NCO1,tplhl$CI1$NCO1);

     if (A == 1'b1 && CI1 == 1'b1 && CI2 == 1'b1 && CS == 1'b1)
       (B *> S) = (tpllh$B$S$A_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1, tphhl$B$S$A_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1);
     if (A == 1'b1 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b1)
       (B *> S) = (tphlh$B$S$A_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1, tplhl$B$S$A_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1);
     if (A == 1'b1 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b0)
       (B *> S) = (tpllh$B$S$A_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0, tphhl$B$S$A_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0);
     if (A == 1'b1 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b1)
       (B *> S) = (tpllh$B$S$A_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1, tphhl$B$S$A_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1);
     if (A == 1'b1 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b0)
       (B *> S) = (tphlh$B$S$A_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0, tplhl$B$S$A_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0);
     if (A == 1'b1 && CI1 == 1'b0 && CI2 == 1'b0 && CS == 1'b0)
       (B *> S) = (tphlh$B$S$A_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0, tplhl$B$S$A_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0);
     if (A == 1'b0 && CI1 == 1'b1 && CI2 == 1'b1 && CS == 1'b1)
       (B *> S) = (tphlh$B$S$A_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1, tplhl$B$S$A_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1);
     if (A == 1'b0 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b1)
       (B *> S) = (tpllh$B$S$A_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1, tphhl$B$S$A_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1);
     if (A == 1'b0 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b0)
       (B *> S) = (tphlh$B$S$A_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0, tplhl$B$S$A_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0);
     if (A == 1'b0 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b1)
       (B *> S) = (tphlh$B$S$A_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1, tplhl$B$S$A_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1);
     if (A == 1'b0 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b0)
       (B *> S) = (tpllh$B$S$A_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0, tphhl$B$S$A_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0);
     if (A == 1'b0 && CI1 == 1'b0 && CI2 == 1'b0 && CS == 1'b0)
       (B *> S) = (tpllh$B$S$A_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0, tphhl$B$S$A_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0);
     ifnone
       (B *> S) = (tpllh$B$S,tplhl$B$S);

     if (A == 1'b1 && CI2 == 1'b0)
       (B *> NCO2) = (tphlh$B$NCO2$A_EQ_1_AN_CI2_EQ_0, tplhl$B$NCO2$A_EQ_1_AN_CI2_EQ_0);
     if (A == 1'b0 && CI2 == 1'b1)
       (B *> NCO2) = (tphlh$B$NCO2$A_EQ_0_AN_CI2_EQ_1, tplhl$B$NCO2$A_EQ_0_AN_CI2_EQ_1);
     ifnone
       (B *> NCO2) = (tphlh$B$NCO2,tplhl$B$NCO2);

     if (A == 1'b1 && CI1 == 1'b0)
       (B *> NCO1) = (tphlh$B$NCO1$A_EQ_1_AN_CI1_EQ_0, tplhl$B$NCO1$A_EQ_1_AN_CI1_EQ_0);
     if (A == 1'b0 && CI1 == 1'b1)
       (B *> NCO1) = (tphlh$B$NCO1$A_EQ_0_AN_CI1_EQ_1, tplhl$B$NCO1$A_EQ_0_AN_CI1_EQ_1);
     ifnone
       (B *> NCO1) = (tphlh$B$NCO1,tplhl$B$NCO1);

     if (B == 1'b1 && CI1 == 1'b1 && CI2 == 1'b1 && CS == 1'b1)
       (A *> S) = (tpllh$A$S$B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1, tphhl$A$S$B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1);
     if (B == 1'b1 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b1)
       (A *> S) = (tphlh$A$S$B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1, tplhl$A$S$B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1);
     if (B == 1'b1 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b0)
       (A *> S) = (tpllh$A$S$B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0, tphhl$A$S$B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0);
     if (B == 1'b1 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b1)
       (A *> S) = (tpllh$A$S$B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1, tphhl$A$S$B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1);
     if (B == 1'b1 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b0)
       (A *> S) = (tphlh$A$S$B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0, tplhl$A$S$B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0);
     if (B == 1'b1 && CI1 == 1'b0 && CI2 == 1'b0 && CS == 1'b0)
       (A *> S) = (tphlh$A$S$B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0, tplhl$A$S$B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0);
     if (B == 1'b0 && CI1 == 1'b1 && CI2 == 1'b1 && CS == 1'b1)
       (A *> S) = (tphlh$A$S$B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1, tplhl$A$S$B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1);
     if (B == 1'b0 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b1)
       (A *> S) = (tpllh$A$S$B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1, tphhl$A$S$B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1);
     if (B == 1'b0 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b0)
       (A *> S) = (tphlh$A$S$B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0, tplhl$A$S$B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0);
     if (B == 1'b0 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b1)
       (A *> S) = (tphlh$A$S$B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1, tplhl$A$S$B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1);
     if (B == 1'b0 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b0)
       (A *> S) = (tpllh$A$S$B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0, tphhl$A$S$B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0);
     if (B == 1'b0 && CI1 == 1'b0 && CI2 == 1'b0 && CS == 1'b0)
       (A *> S) = (tpllh$A$S$B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0, tphhl$A$S$B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0);
     ifnone
       (A *> S) = (tpllh$A$S,tplhl$A$S);

     if (B == 1'b1 && CI2 == 1'b0)
       (A *> NCO2) = (tphlh$A$NCO2$B_EQ_1_AN_CI2_EQ_0, tplhl$A$NCO2$B_EQ_1_AN_CI2_EQ_0);
     if (B == 1'b0 && CI2 == 1'b1)
       (A *> NCO2) = (tphlh$A$NCO2$B_EQ_0_AN_CI2_EQ_1, tplhl$A$NCO2$B_EQ_0_AN_CI2_EQ_1);
     ifnone
       (A *> NCO2) = (tphlh$A$NCO2,tplhl$A$NCO2);

     if (B == 1'b1 && CI1 == 1'b0)
       (A *> NCO1) = (tphlh$A$NCO1$B_EQ_1_AN_CI1_EQ_0, tplhl$A$NCO1$B_EQ_1_AN_CI1_EQ_0);
     if (B == 1'b0 && CI1 == 1'b1)
       (A *> NCO1) = (tphlh$A$NCO1$B_EQ_0_AN_CI1_EQ_1, tplhl$A$NCO1$B_EQ_0_AN_CI1_EQ_1);
     ifnone
       (A *> NCO1) = (tphlh$A$NCO1,tplhl$A$NCO1);*/

// path delays
      (posedge A => (S +: S)) = (1.0, 1.0);
      (negedge A => (S -: S)) = (1.0, 1.0);
      if (B == 1'b0 && CI1 == 1'b1) (A -=> NCO1) = (1.0, 1.0);
      if (B == 1'b1 && CI1 == 1'b0) (A -=> NCO1) = (1.0, 1.0);

      if (B == 1'b1 && CI2 == 1'b0) (A -=> NCO2) = (1.0, 1.0);
      if (B == 1'b0 && CI2 == 1'b1) (A -=> NCO2) = (1.0, 1.0);


      if (B == 1'b1 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b1) (A +=> S) = (1.0, 1.0);
      if (B == 1'b1 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b0) (A +=> S) = (1.0, 1.0);
      if (B == 1'b1 && CI1 == 1'b1 && CI2 == 1'b1 && CS == 1'b1) (A +=> S) = (1.0, 1.0);
      if (B == 1'b0 && CI1 == 1'b0 && CI2 == 1'b0 && CS == 1'b0) (A +=> S) = (1.0, 1.0);
      if (B == 1'b0 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b1) (A +=> S) = (1.0, 1.0);
      if (B == 1'b0 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b0) (A +=> S) = (1.0, 1.0);
   

      if (B == 1'b0 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b1) (A -=> S) = (1.0, 1.0);
      if (B == 1'b0 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b0) (A -=> S) = (1.0, 1.0);
      if (B == 1'b1 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b1) (A -=> S) = (1.0, 1.0);
      if (B == 1'b1 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b0) (A -=> S) = (1.0, 1.0);
      if (B == 1'b1 && CI1 == 1'b0 && CI2 == 1'b0 && CS == 1'b0) (A -=> S) = (1.0, 1.0);
      if (B == 1'b0 && CI1 == 1'b1 && CI2 == 1'b1 && CS == 1'b1) (A -=> S) = (1.0, 1.0);

      (posedge B => (S +: S)) = (1.0, 1.0);
      (negedge B => (S -: S)) = (1.0, 1.0);
      if (A == 1'b1 && CI1 == 1'b0) (B -=> NCO1) = (1.0, 1.0);
      if (A == 1'b0 && CI1 == 1'b1) (B -=> NCO1) = (1.0, 1.0);
  
      if (A == 1'b1 && CI2 == 1'b0) (B -=> NCO2) = (1.0, 1.0);
      if (A == 1'b0 && CI2 == 1'b1) (B -=> NCO2) = (1.0, 1.0);
  

      if (A == 1'b1 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b1) (B +=> S) = (1.0, 1.0);
      if (A == 1'b1 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b0) (B +=> S) = (1.0, 1.0);
      if (A == 1'b1 && CI1 == 1'b1 && CI2 == 1'b1 && CS == 1'b1) (B +=> S) = (1.0, 1.0);
      if (A == 1'b0 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b1) (B +=> S) = (1.0, 1.0);
      if (A == 1'b0 && CI1 == 1'b0 && CI2 == 1'b0 && CS == 1'b0) (B +=> S) = (1.0, 1.0);
      if (A == 1'b0 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b0) (B +=> S) = (1.0, 1.0);
   

      if (A == 1'b0 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b1) (B -=> S) = (1.0, 1.0);
      if (A == 1'b0 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b0) (B -=> S) = (1.0, 1.0);
      if (A == 1'b1 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b1) (B -=> S) = (1.0, 1.0);
      if (A == 1'b1 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b0) (B -=> S) = (1.0, 1.0);
      if (A == 1'b1 && CI1 == 1'b0 && CI2 == 1'b0 && CS == 1'b0) (B -=> S) = (1.0, 1.0);
      if (A == 1'b0 && CI1 == 1'b1 && CI2 == 1'b1 && CS == 1'b1) (B -=> S) = (1.0, 1.0);


      (posedge CI1 => (S +: S)) = (1.0, 1.0);
      (negedge CI1 => (S -: S)) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1) (CI1 -=> NCO1) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0) (CI1 -=> NCO1) = (1.0, 1.0);

      
      if (A == 1'b1 && B == 1'b1 && CI2 == 1'b1 && CS == 1'b0) (CI1 +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b0 && CI2 == 1'b0 && CS == 1'b0) (CI1 +=> S) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0 && CI2 == 1'b0 && CS == 1'b0) (CI1 -=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1 && CI2 == 1'b0 && CS == 1'b0) (CI1 -=> S) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0 && CI2 == 1'b1 && CS == 1'b0) (CI1 -=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1 && CI2 == 1'b1 && CS == 1'b0) (CI1 -=> S) = (1.0, 1.0);
   

      (posedge CI2 => (S +: S)) = (1.0, 1.0);
      (negedge CI2 => (S -: S)) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1) (CI2 -=> NCO2) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0) (CI2 -=> NCO2) = (1.0, 1.0);

      if (A == 1'b1 && B == 1'b1 && CI1 == 1'b1 && CS == 1'b1) (CI2 +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b0 && CI1 == 1'b0 && CS == 1'b1) (CI2 +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1 && CI1 == 1'b0 && CS == 1'b1) (CI2 -=> S) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0 && CI1 == 1'b0 && CS == 1'b1) (CI2 -=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1 && CI1 == 1'b1 && CS == 1'b1) (CI2 -=> S) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0 && CI1 == 1'b1 && CS == 1'b1) (CI2 -=> S) = (1.0, 1.0);

      (posedge CS => (S +: S)) = (1.0, 1.0);
      (negedge CS => (S -: S)) = (1.0, 1.0);

      if (A == 1'b1 && B == 1'b1 && CI1 == 1'b0 && CI2 == 1'b1) (CS +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b0 && CI1 == 1'b0 && CI2 == 1'b1) (CS +=> S) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b1 && CI1 == 1'b1 && CI2 == 1'b0) (CS -=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b0 && CI1 == 1'b1 && CI2 == 1'b0) (CS -=> S) = (1.0, 1.0);
     
   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_FA04D2 (NCO1, NCO2, S, A, B, CI1, CI2, CS);
input  A ;
input  B ;
input  CI1 ;
input  CI2 ;
input  CS ;
output NCO1 ;
output NCO2 ;
output S ;

   and (I0_out, A, B);
   and (I1_out, B, CI1);
   and (I3_out, CI1, A);
   or  (I4_out, I0_out, I1_out, I3_out);
   not (NCO1, I4_out);
   and (I6_out, A, B);
   and (I7_out, B, CI2);
   and (I9_out, CI2, A);
   or  (I10_out, I6_out, I7_out, I9_out);
   not (NCO2, I10_out);
   udp_mux2 (I12_out, CI1, CI2, CS);
   xor (I13_out, I12_out, A);
   xor (S, I13_out, B);

   specify
     // delay parameters
   /*  specparam
       tpllh$A$S = 1.0,
       tplhl$A$S = 1.0,
       tphlh$A$S = 1.0,
       tphhl$A$S = 1.0,
       tplhl$A$NCO2 = 1.0,
       tphlh$A$NCO2 = 1.0,
       tplhl$A$NCO1 = 1.0,
       tphlh$A$NCO1 = 1.0,
       tpllh$B$S = 1.0,
       tplhl$B$S = 1.0,
       tphlh$B$S = 1.0,
       tphhl$B$S = 1.0,
       tplhl$B$NCO2 = 1.0,
       tphlh$B$NCO2 = 1.0,
       tplhl$B$NCO1 = 1.0,
       tphlh$B$NCO1 = 1.0,
       tpllh$CI1$S = 1.0,
       tplhl$CI1$S = 1.0,
       tphlh$CI1$S = 1.0,
       tphhl$CI1$S = 1.0,
       tplhl$CI1$NCO1 = 1.0,
       tphlh$CI1$NCO1 = 1.0,
       tpllh$CI2$S = 1.0,
       tplhl$CI2$S = 1.0,
       tphlh$CI2$S = 1.0,
       tphhl$CI2$S = 1.0,
       tplhl$CI2$NCO2 = 1.0,
       tphlh$CI2$NCO2 = 1.0,
       tpllh$CS$S = 1.0,
       tplhl$CS$S = 1.0,
       tphlh$CS$S = 1.0,
       tphhl$CS$S = 1.0,
       tpllh$A$S$B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tphhl$A$S$B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tpllh$A$S$B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tphhl$A$S$B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tpllh$A$S$B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tphhl$A$S$B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tpllh$A$S$B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tphhl$A$S$B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tpllh$A$S$B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1 = 1.0,
       tphhl$A$S$B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1 = 1.0,
       tpllh$A$S$B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tphhl$A$S$B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tplhl$A$S$B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tphlh$A$S$B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tplhl$A$S$B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1 = 1.0,
       tphlh$A$S$B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1 = 1.0,
       tplhl$A$S$B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tphlh$A$S$B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tplhl$A$S$B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tphlh$A$S$B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tplhl$A$S$B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tphlh$A$S$B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tplhl$A$S$B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tphlh$A$S$B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tplhl$A$NCO2$B_EQ_1_AN_CI2_EQ_0 = 1.0,
       tphlh$A$NCO2$B_EQ_1_AN_CI2_EQ_0 = 1.0,
       tplhl$A$NCO2$B_EQ_0_AN_CI2_EQ_1 = 1.0,
       tphlh$A$NCO2$B_EQ_0_AN_CI2_EQ_1 = 1.0,
       tplhl$A$NCO1$B_EQ_1_AN_CI1_EQ_0 = 1.0,
       tphlh$A$NCO1$B_EQ_1_AN_CI1_EQ_0 = 1.0,
       tplhl$A$NCO1$B_EQ_0_AN_CI1_EQ_1 = 1.0,
       tphlh$A$NCO1$B_EQ_0_AN_CI1_EQ_1 = 1.0,
       tpllh$B$S$A_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tphhl$B$S$A_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tpllh$B$S$A_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tphhl$B$S$A_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tpllh$B$S$A_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tphhl$B$S$A_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tpllh$B$S$A_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tphhl$B$S$A_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tpllh$B$S$A_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1 = 1.0,
       tphhl$B$S$A_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1 = 1.0,
       tpllh$B$S$A_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tphhl$B$S$A_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tplhl$B$S$A_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tphlh$B$S$A_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tplhl$B$S$A_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tphlh$B$S$A_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tplhl$B$S$A_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1 = 1.0,
       tphlh$B$S$A_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1 = 1.0,
       tplhl$B$S$A_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tphlh$B$S$A_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tplhl$B$S$A_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tphlh$B$S$A_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tplhl$B$S$A_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tphlh$B$S$A_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tplhl$B$NCO2$A_EQ_1_AN_CI2_EQ_0 = 1.0,
       tphlh$B$NCO2$A_EQ_1_AN_CI2_EQ_0 = 1.0,
       tplhl$B$NCO2$A_EQ_0_AN_CI2_EQ_1 = 1.0,
       tphlh$B$NCO2$A_EQ_0_AN_CI2_EQ_1 = 1.0,
       tplhl$B$NCO1$A_EQ_1_AN_CI1_EQ_0 = 1.0,
       tphlh$B$NCO1$A_EQ_1_AN_CI1_EQ_0 = 1.0,
       tplhl$B$NCO1$A_EQ_0_AN_CI1_EQ_1 = 1.0,
       tphlh$B$NCO1$A_EQ_0_AN_CI1_EQ_1 = 1.0,
       tpllh$CI1$S$A_EQ_1_AN_B_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tphhl$CI1$S$A_EQ_1_AN_B_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tpllh$CI1$S$A_EQ_0_AN_B_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tphhl$CI1$S$A_EQ_0_AN_B_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tplhl$CI1$S$A_EQ_1_AN_B_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tphlh$CI1$S$A_EQ_1_AN_B_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tplhl$CI1$S$A_EQ_0_AN_B_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tphlh$CI1$S$A_EQ_0_AN_B_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tplhl$CI1$S$A_EQ_1_AN_B_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tphlh$CI1$S$A_EQ_1_AN_B_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tplhl$CI1$S$A_EQ_0_AN_B_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tphlh$CI1$S$A_EQ_0_AN_B_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tplhl$CI1$NCO1$A_EQ_0_AN_B_EQ_1 = 1.0,
       tphlh$CI1$NCO1$A_EQ_0_AN_B_EQ_1 = 1.0,
       tplhl$CI1$NCO1$A_EQ_1_AN_B_EQ_0 = 1.0,
       tphlh$CI1$NCO1$A_EQ_1_AN_B_EQ_0 = 1.0,
       tpllh$CI2$S$A_EQ_1_AN_B_EQ_1_AN_CI1_EQ_1_AN_CS_EQ_1 = 1.0,
       tphhl$CI2$S$A_EQ_1_AN_B_EQ_1_AN_CI1_EQ_1_AN_CS_EQ_1 = 1.0,
       tpllh$CI2$S$A_EQ_0_AN_B_EQ_0_AN_CI1_EQ_0_AN_CS_EQ_1 = 1.0,
       tphhl$CI2$S$A_EQ_0_AN_B_EQ_0_AN_CI1_EQ_0_AN_CS_EQ_1 = 1.0,
       tplhl$CI2$S$A_EQ_1_AN_B_EQ_0_AN_CI1_EQ_0_AN_CS_EQ_1 = 1.0,
       tphlh$CI2$S$A_EQ_1_AN_B_EQ_0_AN_CI1_EQ_0_AN_CS_EQ_1 = 1.0,
       tplhl$CI2$S$A_EQ_0_AN_B_EQ_1_AN_CI1_EQ_0_AN_CS_EQ_1 = 1.0,
       tphlh$CI2$S$A_EQ_0_AN_B_EQ_1_AN_CI1_EQ_0_AN_CS_EQ_1 = 1.0,
       tplhl$CI2$S$A_EQ_1_AN_B_EQ_0_AN_CI1_EQ_1_AN_CS_EQ_1 = 1.0,
       tphlh$CI2$S$A_EQ_1_AN_B_EQ_0_AN_CI1_EQ_1_AN_CS_EQ_1 = 1.0,
       tplhl$CI2$S$A_EQ_0_AN_B_EQ_1_AN_CI1_EQ_1_AN_CS_EQ_1 = 1.0,
       tphlh$CI2$S$A_EQ_0_AN_B_EQ_1_AN_CI1_EQ_1_AN_CS_EQ_1 = 1.0,
       tplhl$CI2$NCO2$A_EQ_0_AN_B_EQ_1 = 1.0,
       tphlh$CI2$NCO2$A_EQ_0_AN_B_EQ_1 = 1.0,
       tplhl$CI2$NCO2$A_EQ_1_AN_B_EQ_0 = 1.0,
       tphlh$CI2$NCO2$A_EQ_1_AN_B_EQ_0 = 1.0,
       tpllh$CS$S$A_EQ_0_AN_B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1 = 1.0,
       tphhl$CS$S$A_EQ_0_AN_B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1 = 1.0,
       tpllh$CS$S$A_EQ_1_AN_B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1 = 1.0,
       tphhl$CS$S$A_EQ_1_AN_B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1 = 1.0,
       tplhl$CS$S$A_EQ_1_AN_B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0 = 1.0,
       tphlh$CS$S$A_EQ_1_AN_B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0 = 1.0,
       tplhl$CS$S$A_EQ_0_AN_B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0 = 1.0,
       tphlh$CS$S$A_EQ_0_AN_B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0 = 1.0;

     // path delays
     if (A == 1'b1 && B == 1'b1 && CI1 == 1'b1 && CI2 == 1'b0)
       (CS *> S) = (tphlh$CS$S$A_EQ_1_AN_B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0, tplhl$CS$S$A_EQ_1_AN_B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0);
     if (A == 1'b1 && B == 1'b1 && CI1 == 1'b0 && CI2 == 1'b1)
       (CS *> S) = (tpllh$CS$S$A_EQ_1_AN_B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1, tphhl$CS$S$A_EQ_1_AN_B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1);
     if (A == 1'b0 && B == 1'b0 && CI1 == 1'b1 && CI2 == 1'b0)
       (CS *> S) = (tphlh$CS$S$A_EQ_0_AN_B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0, tplhl$CS$S$A_EQ_0_AN_B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0);
     if (A == 1'b0 && B == 1'b0 && CI1 == 1'b0 && CI2 == 1'b1)
       (CS *> S) = (tpllh$CS$S$A_EQ_0_AN_B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1, tphhl$CS$S$A_EQ_0_AN_B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1);
     ifnone
       (CS *> S) = (tpllh$CS$S,tplhl$CS$S);

     if (A == 1'b1 && B == 1'b1 && CI1 == 1'b1 && CS == 1'b1)
       (CI2 *> S) = (tpllh$CI2$S$A_EQ_1_AN_B_EQ_1_AN_CI1_EQ_1_AN_CS_EQ_1, tphhl$CI2$S$A_EQ_1_AN_B_EQ_1_AN_CI1_EQ_1_AN_CS_EQ_1);
     if (A == 1'b1 && B == 1'b0 && CI1 == 1'b1 && CS == 1'b1)
       (CI2 *> S) = (tphlh$CI2$S$A_EQ_1_AN_B_EQ_0_AN_CI1_EQ_1_AN_CS_EQ_1, tplhl$CI2$S$A_EQ_1_AN_B_EQ_0_AN_CI1_EQ_1_AN_CS_EQ_1);
     if (A == 1'b1 && B == 1'b0 && CI1 == 1'b0 && CS == 1'b1)
       (CI2 *> S) = (tphlh$CI2$S$A_EQ_1_AN_B_EQ_0_AN_CI1_EQ_0_AN_CS_EQ_1, tplhl$CI2$S$A_EQ_1_AN_B_EQ_0_AN_CI1_EQ_0_AN_CS_EQ_1);
     if (A == 1'b0 && B == 1'b1 && CI1 == 1'b1 && CS == 1'b1)
       (CI2 *> S) = (tphlh$CI2$S$A_EQ_0_AN_B_EQ_1_AN_CI1_EQ_1_AN_CS_EQ_1, tplhl$CI2$S$A_EQ_0_AN_B_EQ_1_AN_CI1_EQ_1_AN_CS_EQ_1);
     if (A == 1'b0 && B == 1'b1 && CI1 == 1'b0 && CS == 1'b1)
       (CI2 *> S) = (tphlh$CI2$S$A_EQ_0_AN_B_EQ_1_AN_CI1_EQ_0_AN_CS_EQ_1, tplhl$CI2$S$A_EQ_0_AN_B_EQ_1_AN_CI1_EQ_0_AN_CS_EQ_1);
     if (A == 1'b0 && B == 1'b0 && CI1 == 1'b0 && CS == 1'b1)
       (CI2 *> S) = (tpllh$CI2$S$A_EQ_0_AN_B_EQ_0_AN_CI1_EQ_0_AN_CS_EQ_1, tphhl$CI2$S$A_EQ_0_AN_B_EQ_0_AN_CI1_EQ_0_AN_CS_EQ_1);
     ifnone
       (CI2 *> S) = (tpllh$CI2$S,tplhl$CI2$S);

     if (A == 1'b1 && B == 1'b0)
       (CI2 *> NCO2) = (tphlh$CI2$NCO2$A_EQ_1_AN_B_EQ_0, tplhl$CI2$NCO2$A_EQ_1_AN_B_EQ_0);
     if (A == 1'b0 && B == 1'b1)
       (CI2 *> NCO2) = (tphlh$CI2$NCO2$A_EQ_0_AN_B_EQ_1, tplhl$CI2$NCO2$A_EQ_0_AN_B_EQ_1);
     ifnone
       (CI2 *> NCO2) = (tphlh$CI2$NCO2,tplhl$CI2$NCO2);

     if (A == 1'b1 && B == 1'b1 && CI2 == 1'b1 && CS == 1'b0)
       (CI1 *> S) = (tpllh$CI1$S$A_EQ_1_AN_B_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_0, tphhl$CI1$S$A_EQ_1_AN_B_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_0);
     if (A == 1'b1 && B == 1'b0 && CI2 == 1'b1 && CS == 1'b0)
       (CI1 *> S) = (tphlh$CI1$S$A_EQ_1_AN_B_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0, tplhl$CI1$S$A_EQ_1_AN_B_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0);
     if (A == 1'b1 && B == 1'b0 && CI2 == 1'b0 && CS == 1'b0)
       (CI1 *> S) = (tphlh$CI1$S$A_EQ_1_AN_B_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0, tplhl$CI1$S$A_EQ_1_AN_B_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0);
     if (A == 1'b0 && B == 1'b1 && CI2 == 1'b1 && CS == 1'b0)
       (CI1 *> S) = (tphlh$CI1$S$A_EQ_0_AN_B_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_0, tplhl$CI1$S$A_EQ_0_AN_B_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_0);
     if (A == 1'b0 && B == 1'b1 && CI2 == 1'b0 && CS == 1'b0)
       (CI1 *> S) = (tphlh$CI1$S$A_EQ_0_AN_B_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0, tplhl$CI1$S$A_EQ_0_AN_B_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0);
     if (A == 1'b0 && B == 1'b0 && CI2 == 1'b0 && CS == 1'b0)
       (CI1 *> S) = (tpllh$CI1$S$A_EQ_0_AN_B_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0, tphhl$CI1$S$A_EQ_0_AN_B_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0);
     ifnone
       (CI1 *> S) = (tpllh$CI1$S,tplhl$CI1$S);

     if (A == 1'b1 && B == 1'b0)
       (CI1 *> NCO1) = (tphlh$CI1$NCO1$A_EQ_1_AN_B_EQ_0, tplhl$CI1$NCO1$A_EQ_1_AN_B_EQ_0);
     if (A == 1'b0 && B == 1'b1)
       (CI1 *> NCO1) = (tphlh$CI1$NCO1$A_EQ_0_AN_B_EQ_1, tplhl$CI1$NCO1$A_EQ_0_AN_B_EQ_1);
     ifnone
       (CI1 *> NCO1) = (tphlh$CI1$NCO1,tplhl$CI1$NCO1);

     if (A == 1'b1 && CI1 == 1'b1 && CI2 == 1'b1 && CS == 1'b1)
       (B *> S) = (tpllh$B$S$A_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1, tphhl$B$S$A_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1);
     if (A == 1'b1 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b1)
       (B *> S) = (tphlh$B$S$A_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1, tplhl$B$S$A_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1);
     if (A == 1'b1 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b0)
       (B *> S) = (tpllh$B$S$A_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0, tphhl$B$S$A_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0);
     if (A == 1'b1 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b1)
       (B *> S) = (tpllh$B$S$A_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1, tphhl$B$S$A_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1);
     if (A == 1'b1 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b0)
       (B *> S) = (tphlh$B$S$A_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0, tplhl$B$S$A_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0);
     if (A == 1'b1 && CI1 == 1'b0 && CI2 == 1'b0 && CS == 1'b0)
       (B *> S) = (tphlh$B$S$A_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0, tplhl$B$S$A_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0);
     if (A == 1'b0 && CI1 == 1'b1 && CI2 == 1'b1 && CS == 1'b1)
       (B *> S) = (tphlh$B$S$A_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1, tplhl$B$S$A_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1);
     if (A == 1'b0 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b1)
       (B *> S) = (tpllh$B$S$A_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1, tphhl$B$S$A_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1);
     if (A == 1'b0 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b0)
       (B *> S) = (tphlh$B$S$A_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0, tplhl$B$S$A_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0);
     if (A == 1'b0 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b1)
       (B *> S) = (tphlh$B$S$A_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1, tplhl$B$S$A_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1);
     if (A == 1'b0 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b0)
       (B *> S) = (tpllh$B$S$A_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0, tphhl$B$S$A_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0);
     if (A == 1'b0 && CI1 == 1'b0 && CI2 == 1'b0 && CS == 1'b0)
       (B *> S) = (tpllh$B$S$A_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0, tphhl$B$S$A_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0);
     ifnone
       (B *> S) = (tpllh$B$S,tplhl$B$S);

     if (A == 1'b1 && CI2 == 1'b0)
       (B *> NCO2) = (tphlh$B$NCO2$A_EQ_1_AN_CI2_EQ_0, tplhl$B$NCO2$A_EQ_1_AN_CI2_EQ_0);
     if (A == 1'b0 && CI2 == 1'b1)
       (B *> NCO2) = (tphlh$B$NCO2$A_EQ_0_AN_CI2_EQ_1, tplhl$B$NCO2$A_EQ_0_AN_CI2_EQ_1);
     ifnone
       (B *> NCO2) = (tphlh$B$NCO2,tplhl$B$NCO2);

     if (A == 1'b1 && CI1 == 1'b0)
       (B *> NCO1) = (tphlh$B$NCO1$A_EQ_1_AN_CI1_EQ_0, tplhl$B$NCO1$A_EQ_1_AN_CI1_EQ_0);
     if (A == 1'b0 && CI1 == 1'b1)
       (B *> NCO1) = (tphlh$B$NCO1$A_EQ_0_AN_CI1_EQ_1, tplhl$B$NCO1$A_EQ_0_AN_CI1_EQ_1);
     ifnone
       (B *> NCO1) = (tphlh$B$NCO1,tplhl$B$NCO1);

     if (B == 1'b1 && CI1 == 1'b1 && CI2 == 1'b1 && CS == 1'b1)
       (A *> S) = (tpllh$A$S$B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1, tphhl$A$S$B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1);
     if (B == 1'b1 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b1)
       (A *> S) = (tphlh$A$S$B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1, tplhl$A$S$B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1);
     if (B == 1'b1 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b0)
       (A *> S) = (tpllh$A$S$B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0, tphhl$A$S$B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0);
     if (B == 1'b1 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b1)
       (A *> S) = (tpllh$A$S$B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1, tphhl$A$S$B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1);
     if (B == 1'b1 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b0)
       (A *> S) = (tphlh$A$S$B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0, tplhl$A$S$B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0);
     if (B == 1'b1 && CI1 == 1'b0 && CI2 == 1'b0 && CS == 1'b0)
       (A *> S) = (tphlh$A$S$B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0, tplhl$A$S$B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0);
     if (B == 1'b0 && CI1 == 1'b1 && CI2 == 1'b1 && CS == 1'b1)
       (A *> S) = (tphlh$A$S$B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1, tplhl$A$S$B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1);
     if (B == 1'b0 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b1)
       (A *> S) = (tpllh$A$S$B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1, tphhl$A$S$B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1);
     if (B == 1'b0 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b0)
       (A *> S) = (tphlh$A$S$B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0, tplhl$A$S$B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0);
     if (B == 1'b0 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b1)
       (A *> S) = (tphlh$A$S$B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1, tplhl$A$S$B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1);
     if (B == 1'b0 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b0)
       (A *> S) = (tpllh$A$S$B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0, tphhl$A$S$B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0);
     if (B == 1'b0 && CI1 == 1'b0 && CI2 == 1'b0 && CS == 1'b0)
       (A *> S) = (tpllh$A$S$B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0, tphhl$A$S$B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0);
     ifnone
       (A *> S) = (tpllh$A$S,tplhl$A$S);

     if (B == 1'b1 && CI2 == 1'b0)
       (A *> NCO2) = (tphlh$A$NCO2$B_EQ_1_AN_CI2_EQ_0, tplhl$A$NCO2$B_EQ_1_AN_CI2_EQ_0);
     if (B == 1'b0 && CI2 == 1'b1)
       (A *> NCO2) = (tphlh$A$NCO2$B_EQ_0_AN_CI2_EQ_1, tplhl$A$NCO2$B_EQ_0_AN_CI2_EQ_1);
     ifnone
       (A *> NCO2) = (tphlh$A$NCO2,tplhl$A$NCO2);

     if (B == 1'b1 && CI1 == 1'b0)
       (A *> NCO1) = (tphlh$A$NCO1$B_EQ_1_AN_CI1_EQ_0, tplhl$A$NCO1$B_EQ_1_AN_CI1_EQ_0);
     if (B == 1'b0 && CI1 == 1'b1)
       (A *> NCO1) = (tphlh$A$NCO1$B_EQ_0_AN_CI1_EQ_1, tplhl$A$NCO1$B_EQ_0_AN_CI1_EQ_1);
     ifnone
       (A *> NCO1) = (tphlh$A$NCO1,tplhl$A$NCO1);*/

// path delays
      (posedge A => (S +: S)) = (1.0, 1.0);
      (negedge A => (S -: S)) = (1.0, 1.0);
      if (B == 1'b0 && CI1 == 1'b1) (A -=> NCO1) = (1.0, 1.0);
      if (B == 1'b1 && CI1 == 1'b0) (A -=> NCO1) = (1.0, 1.0);

      if (B == 1'b1 && CI2 == 1'b0) (A -=> NCO2) = (1.0, 1.0);
      if (B == 1'b0 && CI2 == 1'b1) (A -=> NCO2) = (1.0, 1.0);


      if (B == 1'b1 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b1) (A +=> S) = (1.0, 1.0);
      if (B == 1'b1 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b0) (A +=> S) = (1.0, 1.0);
      if (B == 1'b1 && CI1 == 1'b1 && CI2 == 1'b1 && CS == 1'b1) (A +=> S) = (1.0, 1.0);
      if (B == 1'b0 && CI1 == 1'b0 && CI2 == 1'b0 && CS == 1'b0) (A +=> S) = (1.0, 1.0);
      if (B == 1'b0 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b1) (A +=> S) = (1.0, 1.0);
      if (B == 1'b0 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b0) (A +=> S) = (1.0, 1.0);
   

      if (B == 1'b0 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b1) (A -=> S) = (1.0, 1.0);
      if (B == 1'b0 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b0) (A -=> S) = (1.0, 1.0);
      if (B == 1'b1 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b1) (A -=> S) = (1.0, 1.0);
      if (B == 1'b1 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b0) (A -=> S) = (1.0, 1.0);
      if (B == 1'b1 && CI1 == 1'b0 && CI2 == 1'b0 && CS == 1'b0) (A -=> S) = (1.0, 1.0);
      if (B == 1'b0 && CI1 == 1'b1 && CI2 == 1'b1 && CS == 1'b1) (A -=> S) = (1.0, 1.0);

      (posedge B => (S +: S)) = (1.0, 1.0);
      (negedge B => (S -: S)) = (1.0, 1.0);
      if (A == 1'b1 && CI1 == 1'b0) (B -=> NCO1) = (1.0, 1.0);
      if (A == 1'b0 && CI1 == 1'b1) (B -=> NCO1) = (1.0, 1.0);
  
      if (A == 1'b1 && CI2 == 1'b0) (B -=> NCO2) = (1.0, 1.0);
      if (A == 1'b0 && CI2 == 1'b1) (B -=> NCO2) = (1.0, 1.0);
  

      if (A == 1'b1 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b1) (B +=> S) = (1.0, 1.0);
      if (A == 1'b1 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b0) (B +=> S) = (1.0, 1.0);
      if (A == 1'b1 && CI1 == 1'b1 && CI2 == 1'b1 && CS == 1'b1) (B +=> S) = (1.0, 1.0);
      if (A == 1'b0 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b1) (B +=> S) = (1.0, 1.0);
      if (A == 1'b0 && CI1 == 1'b0 && CI2 == 1'b0 && CS == 1'b0) (B +=> S) = (1.0, 1.0);
      if (A == 1'b0 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b0) (B +=> S) = (1.0, 1.0);
   

      if (A == 1'b0 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b1) (B -=> S) = (1.0, 1.0);
      if (A == 1'b0 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b0) (B -=> S) = (1.0, 1.0);
      if (A == 1'b1 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b1) (B -=> S) = (1.0, 1.0);
      if (A == 1'b1 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b0) (B -=> S) = (1.0, 1.0);
      if (A == 1'b1 && CI1 == 1'b0 && CI2 == 1'b0 && CS == 1'b0) (B -=> S) = (1.0, 1.0);
      if (A == 1'b0 && CI1 == 1'b1 && CI2 == 1'b1 && CS == 1'b1) (B -=> S) = (1.0, 1.0);


      (posedge CI1 => (S +: S)) = (1.0, 1.0);
      (negedge CI1 => (S -: S)) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1) (CI1 -=> NCO1) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0) (CI1 -=> NCO1) = (1.0, 1.0);

      
      if (A == 1'b1 && B == 1'b1 && CI2 == 1'b1 && CS == 1'b0) (CI1 +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b0 && CI2 == 1'b0 && CS == 1'b0) (CI1 +=> S) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0 && CI2 == 1'b0 && CS == 1'b0) (CI1 -=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1 && CI2 == 1'b0 && CS == 1'b0) (CI1 -=> S) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0 && CI2 == 1'b1 && CS == 1'b0) (CI1 -=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1 && CI2 == 1'b1 && CS == 1'b0) (CI1 -=> S) = (1.0, 1.0);
   

      (posedge CI2 => (S +: S)) = (1.0, 1.0);
      (negedge CI2 => (S -: S)) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1) (CI2 -=> NCO2) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0) (CI2 -=> NCO2) = (1.0, 1.0);

      if (A == 1'b1 && B == 1'b1 && CI1 == 1'b1 && CS == 1'b1) (CI2 +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b0 && CI1 == 1'b0 && CS == 1'b1) (CI2 +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1 && CI1 == 1'b0 && CS == 1'b1) (CI2 -=> S) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0 && CI1 == 1'b0 && CS == 1'b1) (CI2 -=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1 && CI1 == 1'b1 && CS == 1'b1) (CI2 -=> S) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0 && CI1 == 1'b1 && CS == 1'b1) (CI2 -=> S) = (1.0, 1.0);

      (posedge CS => (S +: S)) = (1.0, 1.0);
      (negedge CS => (S -: S)) = (1.0, 1.0);

      if (A == 1'b1 && B == 1'b1 && CI1 == 1'b0 && CI2 == 1'b1) (CS +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b0 && CI1 == 1'b0 && CI2 == 1'b1) (CS +=> S) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b1 && CI1 == 1'b1 && CI2 == 1'b0) (CS -=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b0 && CI1 == 1'b1 && CI2 == 1'b0) (CS -=> S) = (1.0, 1.0);
     




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_FA04D4 (NCO1, NCO2, S, A, B, CI1, CI2, CS);
input  A ;
input  B ;
input  CI1 ;
input  CI2 ;
input  CS ;
output NCO1 ;
output NCO2 ;
output S ;

   and (I0_out, A, B);
   and (I1_out, B, CI1);
   and (I3_out, CI1, A);
   or  (I4_out, I0_out, I1_out, I3_out);
   not (NCO1, I4_out);
   and (I6_out, A, B);
   and (I7_out, B, CI2);
   and (I9_out, CI2, A);
   or  (I10_out, I6_out, I7_out, I9_out);
   not (NCO2, I10_out);
   udp_mux2 (I12_out, CI1, CI2, CS);
   xor (I13_out, I12_out, A);
   xor (S, I13_out, B);

   specify
     // delay parameters
  /*   specparam
       tpllh$A$S = 1.0,
       tplhl$A$S = 1.0,
       tphlh$A$S = 1.0,
       tphhl$A$S = 1.0,
       tplhl$A$NCO2 = 1.0,
       tphlh$A$NCO2 = 1.0,
       tplhl$A$NCO1 = 1.0,
       tphlh$A$NCO1 = 1.0,
       tpllh$B$S = 1.0,
       tplhl$B$S = 1.0,
       tphlh$B$S = 1.0,
       tphhl$B$S = 1.0,
       tplhl$B$NCO2 = 1.0,
       tphlh$B$NCO2 = 1.0,
       tplhl$B$NCO1 = 1.0,
       tphlh$B$NCO1 = 1.0,
       tpllh$CI1$S = 1.0,
       tplhl$CI1$S = 1.0,
       tphlh$CI1$S = 1.0,
       tphhl$CI1$S = 1.0,
       tplhl$CI1$NCO1 = 1.0,
       tphlh$CI1$NCO1 = 1.0,
       tpllh$CI2$S = 1.0,
       tplhl$CI2$S = 1.0,
       tphlh$CI2$S = 1.0,
       tphhl$CI2$S = 1.0,
       tplhl$CI2$NCO2 = 1.0,
       tphlh$CI2$NCO2 = 1.0,
       tpllh$CS$S = 1.0,
       tplhl$CS$S = 1.0,
       tphlh$CS$S = 1.0,
       tphhl$CS$S = 1.0,
       tpllh$A$S$B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tphhl$A$S$B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tpllh$A$S$B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tphhl$A$S$B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tpllh$A$S$B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tphhl$A$S$B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tpllh$A$S$B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tphhl$A$S$B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tpllh$A$S$B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1 = 1.0,
       tphhl$A$S$B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1 = 1.0,
       tpllh$A$S$B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tphhl$A$S$B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tplhl$A$S$B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1 = 1.0,
       tphlh$A$S$B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1 = 1.0,
       tplhl$A$S$B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tphlh$A$S$B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tplhl$A$S$B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tphlh$A$S$B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tplhl$A$S$B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tphlh$A$S$B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tplhl$A$S$B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tphlh$A$S$B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tplhl$A$S$B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tphlh$A$S$B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tplhl$A$NCO2$B_EQ_1_AN_CI2_EQ_0 = 1.0,
       tphlh$A$NCO2$B_EQ_1_AN_CI2_EQ_0 = 1.0,
       tplhl$A$NCO2$B_EQ_0_AN_CI2_EQ_1 = 1.0,
       tphlh$A$NCO2$B_EQ_0_AN_CI2_EQ_1 = 1.0,
       tplhl$A$NCO1$B_EQ_1_AN_CI1_EQ_0 = 1.0,
       tphlh$A$NCO1$B_EQ_1_AN_CI1_EQ_0 = 1.0,
       tplhl$A$NCO1$B_EQ_0_AN_CI1_EQ_1 = 1.0,
       tphlh$A$NCO1$B_EQ_0_AN_CI1_EQ_1 = 1.0,
       tpllh$B$S$A_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tphhl$B$S$A_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tpllh$B$S$A_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tphhl$B$S$A_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tpllh$B$S$A_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tphhl$B$S$A_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tpllh$B$S$A_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tphhl$B$S$A_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tpllh$B$S$A_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1 = 1.0,
       tphhl$B$S$A_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1 = 1.0,
       tpllh$B$S$A_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tphhl$B$S$A_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tplhl$B$S$A_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tphlh$B$S$A_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tplhl$B$S$A_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1 = 1.0,
       tphlh$B$S$A_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1 = 1.0,
       tplhl$B$S$A_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tphlh$B$S$A_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tplhl$B$S$A_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tphlh$B$S$A_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tplhl$B$S$A_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tphlh$B$S$A_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tplhl$B$S$A_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tphlh$B$S$A_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1 = 1.0,
       tplhl$B$NCO2$A_EQ_1_AN_CI2_EQ_0 = 1.0,
       tphlh$B$NCO2$A_EQ_1_AN_CI2_EQ_0 = 1.0,
       tplhl$B$NCO2$A_EQ_0_AN_CI2_EQ_1 = 1.0,
       tphlh$B$NCO2$A_EQ_0_AN_CI2_EQ_1 = 1.0,
       tplhl$B$NCO1$A_EQ_1_AN_CI1_EQ_0 = 1.0,
       tphlh$B$NCO1$A_EQ_1_AN_CI1_EQ_0 = 1.0,
       tplhl$B$NCO1$A_EQ_0_AN_CI1_EQ_1 = 1.0,
       tphlh$B$NCO1$A_EQ_0_AN_CI1_EQ_1 = 1.0,
       tpllh$CI1$S$A_EQ_1_AN_B_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tphhl$CI1$S$A_EQ_1_AN_B_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tpllh$CI1$S$A_EQ_0_AN_B_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tphhl$CI1$S$A_EQ_0_AN_B_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tplhl$CI1$S$A_EQ_0_AN_B_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tphlh$CI1$S$A_EQ_0_AN_B_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tplhl$CI1$S$A_EQ_1_AN_B_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tphlh$CI1$S$A_EQ_1_AN_B_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0 = 1.0,
       tplhl$CI1$S$A_EQ_0_AN_B_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tphlh$CI1$S$A_EQ_0_AN_B_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tplhl$CI1$S$A_EQ_1_AN_B_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tphlh$CI1$S$A_EQ_1_AN_B_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0 = 1.0,
       tplhl$CI1$NCO1$A_EQ_0_AN_B_EQ_1 = 1.0,
       tphlh$CI1$NCO1$A_EQ_0_AN_B_EQ_1 = 1.0,
       tplhl$CI1$NCO1$A_EQ_1_AN_B_EQ_0 = 1.0,
       tphlh$CI1$NCO1$A_EQ_1_AN_B_EQ_0 = 1.0,
       tpllh$CI2$S$A_EQ_1_AN_B_EQ_1_AN_CI1_EQ_1_AN_CS_EQ_1 = 1.0,
       tphhl$CI2$S$A_EQ_1_AN_B_EQ_1_AN_CI1_EQ_1_AN_CS_EQ_1 = 1.0,
       tpllh$CI2$S$A_EQ_0_AN_B_EQ_0_AN_CI1_EQ_0_AN_CS_EQ_1 = 1.0,
       tphhl$CI2$S$A_EQ_0_AN_B_EQ_0_AN_CI1_EQ_0_AN_CS_EQ_1 = 1.0,
       tplhl$CI2$S$A_EQ_0_AN_B_EQ_1_AN_CI1_EQ_0_AN_CS_EQ_1 = 1.0,
       tphlh$CI2$S$A_EQ_0_AN_B_EQ_1_AN_CI1_EQ_0_AN_CS_EQ_1 = 1.0,
       tplhl$CI2$S$A_EQ_1_AN_B_EQ_0_AN_CI1_EQ_0_AN_CS_EQ_1 = 1.0,
       tphlh$CI2$S$A_EQ_1_AN_B_EQ_0_AN_CI1_EQ_0_AN_CS_EQ_1 = 1.0,
       tplhl$CI2$S$A_EQ_0_AN_B_EQ_1_AN_CI1_EQ_1_AN_CS_EQ_1 = 1.0,
       tphlh$CI2$S$A_EQ_0_AN_B_EQ_1_AN_CI1_EQ_1_AN_CS_EQ_1 = 1.0,
       tplhl$CI2$S$A_EQ_1_AN_B_EQ_0_AN_CI1_EQ_1_AN_CS_EQ_1 = 1.0,
       tphlh$CI2$S$A_EQ_1_AN_B_EQ_0_AN_CI1_EQ_1_AN_CS_EQ_1 = 1.0,
       tplhl$CI2$NCO2$A_EQ_0_AN_B_EQ_1 = 1.0,
       tphlh$CI2$NCO2$A_EQ_0_AN_B_EQ_1 = 1.0,
       tplhl$CI2$NCO2$A_EQ_1_AN_B_EQ_0 = 1.0,
       tphlh$CI2$NCO2$A_EQ_1_AN_B_EQ_0 = 1.0,
       tpllh$CS$S$A_EQ_1_AN_B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1 = 1.0,
       tphhl$CS$S$A_EQ_1_AN_B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1 = 1.0,
       tpllh$CS$S$A_EQ_0_AN_B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1 = 1.0,
       tphhl$CS$S$A_EQ_0_AN_B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1 = 1.0,
       tplhl$CS$S$A_EQ_1_AN_B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0 = 1.0,
       tphlh$CS$S$A_EQ_1_AN_B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0 = 1.0,
       tplhl$CS$S$A_EQ_0_AN_B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0 = 1.0,
       tphlh$CS$S$A_EQ_0_AN_B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0 = 1.0;

     // path delays
     if (A == 1'b1 && B == 1'b1 && CI1 == 1'b1 && CI2 == 1'b0)
       (CS *> S) = (tphlh$CS$S$A_EQ_1_AN_B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0, tplhl$CS$S$A_EQ_1_AN_B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0);
     if (A == 1'b1 && B == 1'b1 && CI1 == 1'b0 && CI2 == 1'b1)
       (CS *> S) = (tpllh$CS$S$A_EQ_1_AN_B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1, tphhl$CS$S$A_EQ_1_AN_B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1);
     if (A == 1'b0 && B == 1'b0 && CI1 == 1'b1 && CI2 == 1'b0)
       (CS *> S) = (tphlh$CS$S$A_EQ_0_AN_B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0, tplhl$CS$S$A_EQ_0_AN_B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0);
     if (A == 1'b0 && B == 1'b0 && CI1 == 1'b0 && CI2 == 1'b1)
       (CS *> S) = (tpllh$CS$S$A_EQ_0_AN_B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1, tphhl$CS$S$A_EQ_0_AN_B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1);
     ifnone
       (CS *> S) = (tpllh$CS$S,tplhl$CS$S);

     if (A == 1'b1 && B == 1'b1 && CI1 == 1'b1 && CS == 1'b1)
       (CI2 *> S) = (tpllh$CI2$S$A_EQ_1_AN_B_EQ_1_AN_CI1_EQ_1_AN_CS_EQ_1, tphhl$CI2$S$A_EQ_1_AN_B_EQ_1_AN_CI1_EQ_1_AN_CS_EQ_1);
     if (A == 1'b1 && B == 1'b0 && CI1 == 1'b1 && CS == 1'b1)
       (CI2 *> S) = (tphlh$CI2$S$A_EQ_1_AN_B_EQ_0_AN_CI1_EQ_1_AN_CS_EQ_1, tplhl$CI2$S$A_EQ_1_AN_B_EQ_0_AN_CI1_EQ_1_AN_CS_EQ_1);
     if (A == 1'b1 && B == 1'b0 && CI1 == 1'b0 && CS == 1'b1)
       (CI2 *> S) = (tphlh$CI2$S$A_EQ_1_AN_B_EQ_0_AN_CI1_EQ_0_AN_CS_EQ_1, tplhl$CI2$S$A_EQ_1_AN_B_EQ_0_AN_CI1_EQ_0_AN_CS_EQ_1);
     if (A == 1'b0 && B == 1'b1 && CI1 == 1'b1 && CS == 1'b1)
       (CI2 *> S) = (tphlh$CI2$S$A_EQ_0_AN_B_EQ_1_AN_CI1_EQ_1_AN_CS_EQ_1, tplhl$CI2$S$A_EQ_0_AN_B_EQ_1_AN_CI1_EQ_1_AN_CS_EQ_1);
     if (A == 1'b0 && B == 1'b1 && CI1 == 1'b0 && CS == 1'b1)
       (CI2 *> S) = (tphlh$CI2$S$A_EQ_0_AN_B_EQ_1_AN_CI1_EQ_0_AN_CS_EQ_1, tplhl$CI2$S$A_EQ_0_AN_B_EQ_1_AN_CI1_EQ_0_AN_CS_EQ_1);
     if (A == 1'b0 && B == 1'b0 && CI1 == 1'b0 && CS == 1'b1)
       (CI2 *> S) = (tpllh$CI2$S$A_EQ_0_AN_B_EQ_0_AN_CI1_EQ_0_AN_CS_EQ_1, tphhl$CI2$S$A_EQ_0_AN_B_EQ_0_AN_CI1_EQ_0_AN_CS_EQ_1);
     ifnone
       (CI2 *> S) = (tpllh$CI2$S,tplhl$CI2$S);

     if (A == 1'b1 && B == 1'b0)
       (CI2 *> NCO2) = (tphlh$CI2$NCO2$A_EQ_1_AN_B_EQ_0, tplhl$CI2$NCO2$A_EQ_1_AN_B_EQ_0);
     if (A == 1'b0 && B == 1'b1)
       (CI2 *> NCO2) = (tphlh$CI2$NCO2$A_EQ_0_AN_B_EQ_1, tplhl$CI2$NCO2$A_EQ_0_AN_B_EQ_1);
     ifnone
       (CI2 *> NCO2) = (tphlh$CI2$NCO2,tplhl$CI2$NCO2);

     if (A == 1'b1 && B == 1'b1 && CI2 == 1'b1 && CS == 1'b0)
       (CI1 *> S) = (tpllh$CI1$S$A_EQ_1_AN_B_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_0, tphhl$CI1$S$A_EQ_1_AN_B_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_0);
     if (A == 1'b1 && B == 1'b0 && CI2 == 1'b1 && CS == 1'b0)
       (CI1 *> S) = (tphlh$CI1$S$A_EQ_1_AN_B_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0, tplhl$CI1$S$A_EQ_1_AN_B_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0);
     if (A == 1'b1 && B == 1'b0 && CI2 == 1'b0 && CS == 1'b0)
       (CI1 *> S) = (tphlh$CI1$S$A_EQ_1_AN_B_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0, tplhl$CI1$S$A_EQ_1_AN_B_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0);
     if (A == 1'b0 && B == 1'b1 && CI2 == 1'b1 && CS == 1'b0)
       (CI1 *> S) = (tphlh$CI1$S$A_EQ_0_AN_B_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_0, tplhl$CI1$S$A_EQ_0_AN_B_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_0);
     if (A == 1'b0 && B == 1'b1 && CI2 == 1'b0 && CS == 1'b0)
       (CI1 *> S) = (tphlh$CI1$S$A_EQ_0_AN_B_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0, tplhl$CI1$S$A_EQ_0_AN_B_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0);
     if (A == 1'b0 && B == 1'b0 && CI2 == 1'b0 && CS == 1'b0)
       (CI1 *> S) = (tpllh$CI1$S$A_EQ_0_AN_B_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0, tphhl$CI1$S$A_EQ_0_AN_B_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0);
     ifnone
       (CI1 *> S) = (tpllh$CI1$S,tplhl$CI1$S);

     if (A == 1'b1 && B == 1'b0)
       (CI1 *> NCO1) = (tphlh$CI1$NCO1$A_EQ_1_AN_B_EQ_0, tplhl$CI1$NCO1$A_EQ_1_AN_B_EQ_0);
     if (A == 1'b0 && B == 1'b1)
       (CI1 *> NCO1) = (tphlh$CI1$NCO1$A_EQ_0_AN_B_EQ_1, tplhl$CI1$NCO1$A_EQ_0_AN_B_EQ_1);
     ifnone
       (CI1 *> NCO1) = (tphlh$CI1$NCO1,tplhl$CI1$NCO1);

     if (A == 1'b1 && CI1 == 1'b1 && CI2 == 1'b1 && CS == 1'b1)
       (B *> S) = (tpllh$B$S$A_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1, tphhl$B$S$A_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1);
     if (A == 1'b1 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b1)
       (B *> S) = (tphlh$B$S$A_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1, tplhl$B$S$A_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1);
     if (A == 1'b1 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b0)
       (B *> S) = (tpllh$B$S$A_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0, tphhl$B$S$A_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0);
     if (A == 1'b1 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b1)
       (B *> S) = (tpllh$B$S$A_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1, tphhl$B$S$A_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1);
     if (A == 1'b1 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b0)
       (B *> S) = (tphlh$B$S$A_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0, tplhl$B$S$A_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0);
     if (A == 1'b1 && CI1 == 1'b0 && CI2 == 1'b0 && CS == 1'b0)
       (B *> S) = (tphlh$B$S$A_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0, tplhl$B$S$A_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0);
     if (A == 1'b0 && CI1 == 1'b1 && CI2 == 1'b1 && CS == 1'b1)
       (B *> S) = (tphlh$B$S$A_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1, tplhl$B$S$A_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1);
     if (A == 1'b0 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b1)
       (B *> S) = (tpllh$B$S$A_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1, tphhl$B$S$A_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1);
     if (A == 1'b0 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b0)
       (B *> S) = (tphlh$B$S$A_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0, tplhl$B$S$A_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0);
     if (A == 1'b0 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b1)
       (B *> S) = (tphlh$B$S$A_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1, tplhl$B$S$A_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1);
     if (A == 1'b0 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b0)
       (B *> S) = (tpllh$B$S$A_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0, tphhl$B$S$A_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0);
     if (A == 1'b0 && CI1 == 1'b0 && CI2 == 1'b0 && CS == 1'b0)
       (B *> S) = (tpllh$B$S$A_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0, tphhl$B$S$A_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0);
     ifnone
       (B *> S) = (tpllh$B$S,tplhl$B$S);

     if (A == 1'b1 && CI2 == 1'b0)
       (B *> NCO2) = (tphlh$B$NCO2$A_EQ_1_AN_CI2_EQ_0, tplhl$B$NCO2$A_EQ_1_AN_CI2_EQ_0);
     if (A == 1'b0 && CI2 == 1'b1)
       (B *> NCO2) = (tphlh$B$NCO2$A_EQ_0_AN_CI2_EQ_1, tplhl$B$NCO2$A_EQ_0_AN_CI2_EQ_1);
     ifnone
       (B *> NCO2) = (tphlh$B$NCO2,tplhl$B$NCO2);

     if (A == 1'b1 && CI1 == 1'b0)
       (B *> NCO1) = (tphlh$B$NCO1$A_EQ_1_AN_CI1_EQ_0, tplhl$B$NCO1$A_EQ_1_AN_CI1_EQ_0);
     if (A == 1'b0 && CI1 == 1'b1)
       (B *> NCO1) = (tphlh$B$NCO1$A_EQ_0_AN_CI1_EQ_1, tplhl$B$NCO1$A_EQ_0_AN_CI1_EQ_1);
     ifnone
       (B *> NCO1) = (tphlh$B$NCO1,tplhl$B$NCO1);

     if (B == 1'b1 && CI1 == 1'b1 && CI2 == 1'b1 && CS == 1'b1)
       (A *> S) = (tpllh$A$S$B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1, tphhl$A$S$B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1);
     if (B == 1'b1 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b1)
       (A *> S) = (tphlh$A$S$B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1, tplhl$A$S$B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1);
     if (B == 1'b1 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b0)
       (A *> S) = (tpllh$A$S$B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0, tphhl$A$S$B_EQ_1_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0);
     if (B == 1'b1 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b1)
       (A *> S) = (tpllh$A$S$B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1, tphhl$A$S$B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1);
     if (B == 1'b1 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b0)
       (A *> S) = (tphlh$A$S$B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0, tplhl$A$S$B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0);
     if (B == 1'b1 && CI1 == 1'b0 && CI2 == 1'b0 && CS == 1'b0)
       (A *> S) = (tphlh$A$S$B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0, tplhl$A$S$B_EQ_1_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0);
     if (B == 1'b0 && CI1 == 1'b1 && CI2 == 1'b1 && CS == 1'b1)
       (A *> S) = (tphlh$A$S$B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1, tplhl$A$S$B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_1_AN_CS_EQ_1);
     if (B == 1'b0 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b1)
       (A *> S) = (tpllh$A$S$B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1, tphhl$A$S$B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_1);
     if (B == 1'b0 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b0)
       (A *> S) = (tphlh$A$S$B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0, tplhl$A$S$B_EQ_0_AN_CI1_EQ_1_AN_CI2_EQ_0_AN_CS_EQ_0);
     if (B == 1'b0 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b1)
       (A *> S) = (tphlh$A$S$B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1, tplhl$A$S$B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_1);
     if (B == 1'b0 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b0)
       (A *> S) = (tpllh$A$S$B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0, tphhl$A$S$B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_1_AN_CS_EQ_0);
     if (B == 1'b0 && CI1 == 1'b0 && CI2 == 1'b0 && CS == 1'b0)
       (A *> S) = (tpllh$A$S$B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0, tphhl$A$S$B_EQ_0_AN_CI1_EQ_0_AN_CI2_EQ_0_AN_CS_EQ_0);
     ifnone
       (A *> S) = (tpllh$A$S,tplhl$A$S);

     if (B == 1'b1 && CI2 == 1'b0)
       (A *> NCO2) = (tphlh$A$NCO2$B_EQ_1_AN_CI2_EQ_0, tplhl$A$NCO2$B_EQ_1_AN_CI2_EQ_0);
     if (B == 1'b0 && CI2 == 1'b1)
       (A *> NCO2) = (tphlh$A$NCO2$B_EQ_0_AN_CI2_EQ_1, tplhl$A$NCO2$B_EQ_0_AN_CI2_EQ_1);
     ifnone
       (A *> NCO2) = (tphlh$A$NCO2,tplhl$A$NCO2);

     if (B == 1'b1 && CI1 == 1'b0)
       (A *> NCO1) = (tphlh$A$NCO1$B_EQ_1_AN_CI1_EQ_0, tplhl$A$NCO1$B_EQ_1_AN_CI1_EQ_0);
     if (B == 1'b0 && CI1 == 1'b1)
       (A *> NCO1) = (tphlh$A$NCO1$B_EQ_0_AN_CI1_EQ_1, tplhl$A$NCO1$B_EQ_0_AN_CI1_EQ_1);
     ifnone
       (A *> NCO1) = (tphlh$A$NCO1,tplhl$A$NCO1);*/

// path delays
      (posedge A => (S +: S)) = (1.0, 1.0);
      (negedge A => (S -: S)) = (1.0, 1.0);
      if (B == 1'b0 && CI1 == 1'b1) (A -=> NCO1) = (1.0, 1.0);
      if (B == 1'b1 && CI1 == 1'b0) (A -=> NCO1) = (1.0, 1.0);

      if (B == 1'b1 && CI2 == 1'b0) (A -=> NCO2) = (1.0, 1.0);
      if (B == 1'b0 && CI2 == 1'b1) (A -=> NCO2) = (1.0, 1.0);


      if (B == 1'b1 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b1) (A +=> S) = (1.0, 1.0);
      if (B == 1'b1 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b0) (A +=> S) = (1.0, 1.0);
      if (B == 1'b1 && CI1 == 1'b1 && CI2 == 1'b1 && CS == 1'b1) (A +=> S) = (1.0, 1.0);
      if (B == 1'b0 && CI1 == 1'b0 && CI2 == 1'b0 && CS == 1'b0) (A +=> S) = (1.0, 1.0);
      if (B == 1'b0 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b1) (A +=> S) = (1.0, 1.0);
      if (B == 1'b0 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b0) (A +=> S) = (1.0, 1.0);
   

      if (B == 1'b0 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b1) (A -=> S) = (1.0, 1.0);
      if (B == 1'b0 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b0) (A -=> S) = (1.0, 1.0);
      if (B == 1'b1 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b1) (A -=> S) = (1.0, 1.0);
      if (B == 1'b1 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b0) (A -=> S) = (1.0, 1.0);
      if (B == 1'b1 && CI1 == 1'b0 && CI2 == 1'b0 && CS == 1'b0) (A -=> S) = (1.0, 1.0);
      if (B == 1'b0 && CI1 == 1'b1 && CI2 == 1'b1 && CS == 1'b1) (A -=> S) = (1.0, 1.0);

      (posedge B => (S +: S)) = (1.0, 1.0);
      (negedge B => (S -: S)) = (1.0, 1.0);
      if (A == 1'b1 && CI1 == 1'b0) (B -=> NCO1) = (1.0, 1.0);
      if (A == 1'b0 && CI1 == 1'b1) (B -=> NCO1) = (1.0, 1.0);
  
      if (A == 1'b1 && CI2 == 1'b0) (B -=> NCO2) = (1.0, 1.0);
      if (A == 1'b0 && CI2 == 1'b1) (B -=> NCO2) = (1.0, 1.0);
  

      if (A == 1'b1 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b1) (B +=> S) = (1.0, 1.0);
      if (A == 1'b1 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b0) (B +=> S) = (1.0, 1.0);
      if (A == 1'b1 && CI1 == 1'b1 && CI2 == 1'b1 && CS == 1'b1) (B +=> S) = (1.0, 1.0);
      if (A == 1'b0 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b1) (B +=> S) = (1.0, 1.0);
      if (A == 1'b0 && CI1 == 1'b0 && CI2 == 1'b0 && CS == 1'b0) (B +=> S) = (1.0, 1.0);
      if (A == 1'b0 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b0) (B +=> S) = (1.0, 1.0);
   

      if (A == 1'b0 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b1) (B -=> S) = (1.0, 1.0);
      if (A == 1'b0 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b0) (B -=> S) = (1.0, 1.0);
      if (A == 1'b1 && CI1 == 1'b1 && CI2 == 1'b0 && CS == 1'b1) (B -=> S) = (1.0, 1.0);
      if (A == 1'b1 && CI1 == 1'b0 && CI2 == 1'b1 && CS == 1'b0) (B -=> S) = (1.0, 1.0);
      if (A == 1'b1 && CI1 == 1'b0 && CI2 == 1'b0 && CS == 1'b0) (B -=> S) = (1.0, 1.0);
      if (A == 1'b0 && CI1 == 1'b1 && CI2 == 1'b1 && CS == 1'b1) (B -=> S) = (1.0, 1.0);


      (posedge CI1 => (S +: S)) = (1.0, 1.0);
      (negedge CI1 => (S -: S)) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1) (CI1 -=> NCO1) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0) (CI1 -=> NCO1) = (1.0, 1.0);

      
      if (A == 1'b1 && B == 1'b1 && CI2 == 1'b1 && CS == 1'b0) (CI1 +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b0 && CI2 == 1'b0 && CS == 1'b0) (CI1 +=> S) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0 && CI2 == 1'b0 && CS == 1'b0) (CI1 -=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1 && CI2 == 1'b0 && CS == 1'b0) (CI1 -=> S) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0 && CI2 == 1'b1 && CS == 1'b0) (CI1 -=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1 && CI2 == 1'b1 && CS == 1'b0) (CI1 -=> S) = (1.0, 1.0);
   

      (posedge CI2 => (S +: S)) = (1.0, 1.0);
      (negedge CI2 => (S -: S)) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1) (CI2 -=> NCO2) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0) (CI2 -=> NCO2) = (1.0, 1.0);

      if (A == 1'b1 && B == 1'b1 && CI1 == 1'b1 && CS == 1'b1) (CI2 +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b0 && CI1 == 1'b0 && CS == 1'b1) (CI2 +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1 && CI1 == 1'b0 && CS == 1'b1) (CI2 -=> S) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0 && CI1 == 1'b0 && CS == 1'b1) (CI2 -=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1 && CI1 == 1'b1 && CS == 1'b1) (CI2 -=> S) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0 && CI1 == 1'b1 && CS == 1'b1) (CI2 -=> S) = (1.0, 1.0);

      (posedge CS => (S +: S)) = (1.0, 1.0);
      (negedge CS => (S -: S)) = (1.0, 1.0);

      if (A == 1'b1 && B == 1'b1 && CI1 == 1'b0 && CI2 == 1'b1) (CS +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b0 && CI1 == 1'b0 && CI2 == 1'b1) (CS +=> S) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b1 && CI1 == 1'b1 && CI2 == 1'b0) (CS -=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b0 && CI1 == 1'b1 && CI2 == 1'b0) (CS -=> S) = (1.0, 1.0);


   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_FA05D1 (CO1, CO2, S, A, B, CS, NCI1, NCI2);
input  A ;
input  B ;
input  CS ;
input  NCI1 ;
input  NCI2 ;
output CO1 ;
output CO2 ;
output S ;

   not (I0_out, NCI1);
   and (I1_out, I0_out, A);
   and (I2_out, A, B);
   not (I4_out, NCI1);
   and (I5_out, B, I4_out);
   or  (CO1, I1_out, I2_out, I5_out);
   not (I7_out, NCI2);
   and (I8_out, I7_out, A);
   and (I9_out, A, B);
   not (I11_out, NCI2);
   and (I12_out, B, I11_out);
   or  (CO2, I8_out, I9_out, I12_out);
   udp_mux2 (I14_out, NCI1, NCI2, CS);
   xor (I15_out, I14_out, A);
   xor (I16_out, I15_out, B);
   not (S, I16_out);

   specify
     // delay parameters
 /*    specparam
       tpllh$A$CO1 = 1.0,
       tphhl$A$CO1 = 1.0,
       tpllh$A$CO2 = 1.0,
       tphhl$A$CO2 = 1.0,
       tpllh$A$S = 1.0,
       tplhl$A$S = 1.0,
       tphlh$A$S = 1.0,
       tphhl$A$S = 1.0,
       tpllh$B$CO1 = 1.0,
       tphhl$B$CO1 = 1.0,
       tpllh$B$CO2 = 1.0,
       tphhl$B$CO2 = 1.0,
       tpllh$B$S = 1.0,
       tplhl$B$S = 1.0,
       tphlh$B$S = 1.0,
       tphhl$B$S = 1.0,
       tpllh$CS$S = 1.0,
       tplhl$CS$S = 1.0,
       tphlh$CS$S = 1.0,
       tphhl$CS$S = 1.0,
       tpllh$NCI1$S = 1.0,
       tplhl$NCI1$S = 1.0,
       tphlh$NCI1$S = 1.0,
       tphhl$NCI1$S = 1.0,
       tplhl$NCI1$CO1 = 1.0,
       tphlh$NCI1$CO1 = 1.0,
       tpllh$NCI2$S = 1.0,
       tplhl$NCI2$S = 1.0,
       tphlh$NCI2$S = 1.0,
       tphhl$NCI2$S = 1.0,
       tplhl$NCI2$CO2 = 1.0,
       tphlh$NCI2$CO2 = 1.0,
       tpllh$A$CO1$B_EQ_1_AN_NCI1_EQ_1 = 1.0,
       tphhl$A$CO1$B_EQ_1_AN_NCI1_EQ_1 = 1.0,
       tpllh$A$CO1$B_EQ_0_AN_NCI1_EQ_0 = 1.0,
       tphhl$A$CO1$B_EQ_0_AN_NCI1_EQ_0 = 1.0,
       tpllh$A$CO2$B_EQ_1_AN_NCI2_EQ_1 = 1.0,
       tphhl$A$CO2$B_EQ_1_AN_NCI2_EQ_1 = 1.0,
       tpllh$A$CO2$B_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tphhl$A$CO2$B_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tpllh$A$S$B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tphhl$A$S$B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tpllh$A$S$B_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tphhl$A$S$B_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tpllh$A$S$B_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tphhl$A$S$B_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tpllh$A$S$B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1 = 1.0,
       tphhl$A$S$B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1 = 1.0,
       tpllh$A$S$B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tphhl$A$S$B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tpllh$A$S$B_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tphhl$A$S$B_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tplhl$A$S$B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tphlh$A$S$B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tplhl$A$S$B_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tphlh$A$S$B_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tplhl$A$S$B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tphlh$A$S$B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tplhl$A$S$B_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tphlh$A$S$B_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tplhl$A$S$B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1 = 1.0,
       tphlh$A$S$B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1 = 1.0,
       tplhl$A$S$B_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tphlh$A$S$B_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tpllh$B$CO1$A_EQ_1_AN_NCI1_EQ_1 = 1.0,
       tphhl$B$CO1$A_EQ_1_AN_NCI1_EQ_1 = 1.0,
       tpllh$B$CO1$A_EQ_0_AN_NCI1_EQ_0 = 1.0,
       tphhl$B$CO1$A_EQ_0_AN_NCI1_EQ_0 = 1.0,
       tpllh$B$CO2$A_EQ_1_AN_NCI2_EQ_1 = 1.0,
       tphhl$B$CO2$A_EQ_1_AN_NCI2_EQ_1 = 1.0,
       tpllh$B$CO2$A_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tphhl$B$CO2$A_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tpllh$B$S$A_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tphhl$B$S$A_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tpllh$B$S$A_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tphhl$B$S$A_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tpllh$B$S$A_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tphhl$B$S$A_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tpllh$B$S$A_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1 = 1.0,
       tphhl$B$S$A_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1 = 1.0,
       tpllh$B$S$A_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tphhl$B$S$A_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tpllh$B$S$A_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tphhl$B$S$A_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tplhl$B$S$A_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tphlh$B$S$A_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tplhl$B$S$A_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tphlh$B$S$A_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tplhl$B$S$A_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tphlh$B$S$A_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tplhl$B$S$A_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tphlh$B$S$A_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tplhl$B$S$A_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1 = 1.0,
       tphlh$B$S$A_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1 = 1.0,
       tplhl$B$S$A_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tphlh$B$S$A_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tpllh$CS$S$A_EQ_1_AN_B_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tphhl$CS$S$A_EQ_1_AN_B_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tpllh$CS$S$A_EQ_0_AN_B_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tphhl$CS$S$A_EQ_0_AN_B_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tplhl$CS$S$A_EQ_1_AN_B_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tphlh$CS$S$A_EQ_1_AN_B_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tplhl$CS$S$A_EQ_0_AN_B_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tphlh$CS$S$A_EQ_0_AN_B_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tpllh$NCI1$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tphhl$NCI1$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tpllh$NCI1$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tphhl$NCI1$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tpllh$NCI1$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tphhl$NCI1$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tpllh$NCI1$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tphhl$NCI1$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tplhl$NCI1$S$A_EQ_0_AN_B_EQ_0_AN_CS_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tphlh$NCI1$S$A_EQ_0_AN_B_EQ_0_AN_CS_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tplhl$NCI1$S$A_EQ_1_AN_B_EQ_1_AN_CS_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tphlh$NCI1$S$A_EQ_1_AN_B_EQ_1_AN_CS_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tplhl$NCI1$CO1$A_EQ_0_AN_B_EQ_1 = 1.0,
       tphlh$NCI1$CO1$A_EQ_0_AN_B_EQ_1 = 1.0,
       tplhl$NCI1$CO1$A_EQ_1_AN_B_EQ_0 = 1.0,
       tphlh$NCI1$CO1$A_EQ_1_AN_B_EQ_0 = 1.0,
       tpllh$NCI2$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1 = 1.0,
       tphhl$NCI2$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1 = 1.0,
       tpllh$NCI2$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1 = 1.0,
       tphhl$NCI2$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1 = 1.0,
       tpllh$NCI2$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0 = 1.0,
       tphhl$NCI2$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0 = 1.0,
       tpllh$NCI2$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_0 = 1.0,
       tphhl$NCI2$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_0 = 1.0,
       tplhl$NCI2$S$A_EQ_0_AN_B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0 = 1.0,
       tphlh$NCI2$S$A_EQ_0_AN_B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0 = 1.0,
       tplhl$NCI2$S$A_EQ_1_AN_B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1 = 1.0,
       tphlh$NCI2$S$A_EQ_1_AN_B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1 = 1.0,
       tplhl$NCI2$CO2$A_EQ_0_AN_B_EQ_1 = 1.0,
       tphlh$NCI2$CO2$A_EQ_0_AN_B_EQ_1 = 1.0,
       tplhl$NCI2$CO2$A_EQ_1_AN_B_EQ_0 = 1.0,
       tphlh$NCI2$CO2$A_EQ_1_AN_B_EQ_0 = 1.0;

     // path delays
     if (A == 1'b1 && B == 1'b1 && CS == 1'b1 && NCI1 == 1'b1)
       (NCI2 *> S) = (tphlh$NCI2$S$A_EQ_1_AN_B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1, tplhl$NCI2$S$A_EQ_1_AN_B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1);
     if (A == 1'b1 && B == 1'b0 && CS == 1'b1 && NCI1 == 1'b1)
       (NCI2 *> S) = (tpllh$NCI2$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1, tphhl$NCI2$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1);
     if (A == 1'b1 && B == 1'b0 && CS == 1'b1 && NCI1 == 1'b0)
       (NCI2 *> S) = (tpllh$NCI2$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0, tphhl$NCI2$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0);
     if (A == 1'b0 && B == 1'b1 && CS == 1'b1 && NCI1 == 1'b1)
       (NCI2 *> S) = (tpllh$NCI2$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1, tphhl$NCI2$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1);
     if (A == 1'b0 && B == 1'b1 && CS == 1'b1 && NCI1 == 1'b0)
       (NCI2 *> S) = (tpllh$NCI2$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_0, tphhl$NCI2$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_0);
     if (A == 1'b0 && B == 1'b0 && CS == 1'b1 && NCI1 == 1'b0)
       (NCI2 *> S) = (tphlh$NCI2$S$A_EQ_0_AN_B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0, tplhl$NCI2$S$A_EQ_0_AN_B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0);
     ifnone
       (NCI2 *> S) = (tpllh$NCI2$S,tplhl$NCI2$S);

     if (A == 1'b1 && B == 1'b0)
       (NCI2 *> CO2) = (tphlh$NCI2$CO2$A_EQ_1_AN_B_EQ_0, tplhl$NCI2$CO2$A_EQ_1_AN_B_EQ_0);
     if (A == 1'b0 && B == 1'b1)
       (NCI2 *> CO2) = (tphlh$NCI2$CO2$A_EQ_0_AN_B_EQ_1, tplhl$NCI2$CO2$A_EQ_0_AN_B_EQ_1);
     ifnone
       (NCI2 *> CO2) = (tphlh$NCI2$CO2,tplhl$NCI2$CO2);

     if (A == 1'b1 && B == 1'b1 && CS == 1'b0 && NCI2 == 1'b1)
       (NCI1 *> S) = (tphlh$NCI1$S$A_EQ_1_AN_B_EQ_1_AN_CS_EQ_0_AN_NCI2_EQ_1, tplhl$NCI1$S$A_EQ_1_AN_B_EQ_1_AN_CS_EQ_0_AN_NCI2_EQ_1);
     if (A == 1'b1 && B == 1'b0 && CS == 1'b0 && NCI2 == 1'b1)
       (NCI1 *> S) = (tpllh$NCI1$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_0_AN_NCI2_EQ_1, tphhl$NCI1$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_0_AN_NCI2_EQ_1);
     if (A == 1'b1 && B == 1'b0 && CS == 1'b0 && NCI2 == 1'b0)
       (NCI1 *> S) = (tpllh$NCI1$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_0_AN_NCI2_EQ_0, tphhl$NCI1$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_0_AN_NCI2_EQ_0);
     if (A == 1'b0 && B == 1'b1 && CS == 1'b0 && NCI2 == 1'b1)
       (NCI1 *> S) = (tpllh$NCI1$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_0_AN_NCI2_EQ_1, tphhl$NCI1$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_0_AN_NCI2_EQ_1);
     if (A == 1'b0 && B == 1'b1 && CS == 1'b0 && NCI2 == 1'b0)
       (NCI1 *> S) = (tpllh$NCI1$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_0_AN_NCI2_EQ_0, tphhl$NCI1$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_0_AN_NCI2_EQ_0);
     if (A == 1'b0 && B == 1'b0 && CS == 1'b0 && NCI2 == 1'b0)
       (NCI1 *> S) = (tphlh$NCI1$S$A_EQ_0_AN_B_EQ_0_AN_CS_EQ_0_AN_NCI2_EQ_0, tplhl$NCI1$S$A_EQ_0_AN_B_EQ_0_AN_CS_EQ_0_AN_NCI2_EQ_0);
     ifnone
       (NCI1 *> S) = (tpllh$NCI1$S,tplhl$NCI1$S);

     if (A == 1'b1 && B == 1'b0)
       (NCI1 *> CO1) = (tphlh$NCI1$CO1$A_EQ_1_AN_B_EQ_0, tplhl$NCI1$CO1$A_EQ_1_AN_B_EQ_0);
     if (A == 1'b0 && B == 1'b1)
       (NCI1 *> CO1) = (tphlh$NCI1$CO1$A_EQ_0_AN_B_EQ_1, tplhl$NCI1$CO1$A_EQ_0_AN_B_EQ_1);
     ifnone
       (NCI1 *> CO1) = (tphlh$NCI1$CO1,tplhl$NCI1$CO1);

     if (A == 1'b1 && B == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b0)
       (CS *> S) = (tpllh$CS$S$A_EQ_1_AN_B_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0, tphhl$CS$S$A_EQ_1_AN_B_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0);
     if (A == 1'b1 && B == 1'b1 && NCI1 == 1'b0 && NCI2 == 1'b1)
       (CS *> S) = (tphlh$CS$S$A_EQ_1_AN_B_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1, tplhl$CS$S$A_EQ_1_AN_B_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1);
     if (A == 1'b0 && B == 1'b0 && NCI1 == 1'b1 && NCI2 == 1'b0)
       (CS *> S) = (tpllh$CS$S$A_EQ_0_AN_B_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0, tphhl$CS$S$A_EQ_0_AN_B_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0);
     if (A == 1'b0 && B == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b1)
       (CS *> S) = (tphlh$CS$S$A_EQ_0_AN_B_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1, tplhl$CS$S$A_EQ_0_AN_B_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1);
     ifnone
       (CS *> S) = (tpllh$CS$S,tplhl$CS$S);

     if (A == 1'b1 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b1)
       (B *> S) = (tphlh$B$S$A_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1, tplhl$B$S$A_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1);
     if (A == 1'b1 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b0)
       (B *> S) = (tpllh$B$S$A_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0, tphhl$B$S$A_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0);
     if (A == 1'b1 && CS == 1'b1 && NCI1 == 1'b0 && NCI2 == 1'b1)
       (B *> S) = (tphlh$B$S$A_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1, tplhl$B$S$A_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1);
     if (A == 1'b1 && CS == 1'b0 && NCI1 == 1'b1 && NCI2 == 1'b0)
       (B *> S) = (tphlh$B$S$A_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0, tplhl$B$S$A_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0);
     if (A == 1'b1 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b1)
       (B *> S) = (tpllh$B$S$A_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1, tphhl$B$S$A_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1);
     if (A == 1'b1 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b0)
       (B *> S) = (tpllh$B$S$A_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0, tphhl$B$S$A_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0);
     if (A == 1'b0 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b1)
       (B *> S) = (tpllh$B$S$A_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1, tphhl$B$S$A_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1);
     if (A == 1'b0 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b0)
       (B *> S) = (tphlh$B$S$A_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0, tplhl$B$S$A_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0);
     if (A == 1'b0 && CS == 1'b1 && NCI1 == 1'b0 && NCI2 == 1'b1)
       (B *> S) = (tpllh$B$S$A_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1, tphhl$B$S$A_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1);
     if (A == 1'b0 && CS == 1'b0 && NCI1 == 1'b1 && NCI2 == 1'b0)
       (B *> S) = (tpllh$B$S$A_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0, tphhl$B$S$A_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0);
     if (A == 1'b0 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b1)
       (B *> S) = (tphlh$B$S$A_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1, tplhl$B$S$A_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1);
     if (A == 1'b0 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b0)
       (B *> S) = (tphlh$B$S$A_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0, tplhl$B$S$A_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0);
     ifnone
       (B *> S) = (tpllh$B$S,tplhl$B$S);

     if (A == 1'b1 && NCI2 == 1'b1)
       (B *> CO2) = (tpllh$B$CO2$A_EQ_1_AN_NCI2_EQ_1, tphhl$B$CO2$A_EQ_1_AN_NCI2_EQ_1);
     if (A == 1'b0 && NCI2 == 1'b0)
       (B *> CO2) = (tpllh$B$CO2$A_EQ_0_AN_NCI2_EQ_0, tphhl$B$CO2$A_EQ_0_AN_NCI2_EQ_0);
     ifnone
       (B *> CO2) = (tpllh$B$CO2,tphhl$B$CO2);

     if (A == 1'b1 && NCI1 == 1'b1)
       (B *> CO1) = (tpllh$B$CO1$A_EQ_1_AN_NCI1_EQ_1, tphhl$B$CO1$A_EQ_1_AN_NCI1_EQ_1);
     if (A == 1'b0 && NCI1 == 1'b0)
       (B *> CO1) = (tpllh$B$CO1$A_EQ_0_AN_NCI1_EQ_0, tphhl$B$CO1$A_EQ_0_AN_NCI1_EQ_0);
     ifnone
       (B *> CO1) = (tpllh$B$CO1,tphhl$B$CO1);

     if (B == 1'b1 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b1)
       (A *> S) = (tphlh$A$S$B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1, tplhl$A$S$B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1);
     if (B == 1'b1 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b0)
       (A *> S) = (tpllh$A$S$B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0, tphhl$A$S$B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0);
     if (B == 1'b1 && CS == 1'b1 && NCI1 == 1'b0 && NCI2 == 1'b1)
       (A *> S) = (tphlh$A$S$B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1, tplhl$A$S$B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1);
     if (B == 1'b1 && CS == 1'b0 && NCI1 == 1'b1 && NCI2 == 1'b0)
       (A *> S) = (tphlh$A$S$B_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0, tplhl$A$S$B_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0);
     if (B == 1'b1 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b1)
       (A *> S) = (tpllh$A$S$B_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1, tphhl$A$S$B_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1);
     if (B == 1'b1 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b0)
       (A *> S) = (tpllh$A$S$B_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0, tphhl$A$S$B_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0);
     if (B == 1'b0 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b1)
       (A *> S) = (tpllh$A$S$B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1, tphhl$A$S$B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1);
     if (B == 1'b0 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b0)
       (A *> S) = (tphlh$A$S$B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0, tplhl$A$S$B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0);
     if (B == 1'b0 && CS == 1'b1 && NCI1 == 1'b0 && NCI2 == 1'b1)
       (A *> S) = (tpllh$A$S$B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1, tphhl$A$S$B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1);
     if (B == 1'b0 && CS == 1'b0 && NCI1 == 1'b1 && NCI2 == 1'b0)
       (A *> S) = (tpllh$A$S$B_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0, tphhl$A$S$B_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0);
     if (B == 1'b0 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b1)
       (A *> S) = (tphlh$A$S$B_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1, tplhl$A$S$B_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1);
     if (B == 1'b0 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b0)
       (A *> S) = (tphlh$A$S$B_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0, tplhl$A$S$B_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0);
     ifnone
       (A *> S) = (tpllh$A$S,tplhl$A$S);

     if (B == 1'b1 && NCI2 == 1'b1)
       (A *> CO2) = (tpllh$A$CO2$B_EQ_1_AN_NCI2_EQ_1, tphhl$A$CO2$B_EQ_1_AN_NCI2_EQ_1);
     if (B == 1'b0 && NCI2 == 1'b0)
       (A *> CO2) = (tpllh$A$CO2$B_EQ_0_AN_NCI2_EQ_0, tphhl$A$CO2$B_EQ_0_AN_NCI2_EQ_0);
     ifnone
       (A *> CO2) = (tpllh$A$CO2,tphhl$A$CO2);

     if (B == 1'b1 && NCI1 == 1'b1)
       (A *> CO1) = (tpllh$A$CO1$B_EQ_1_AN_NCI1_EQ_1, tphhl$A$CO1$B_EQ_1_AN_NCI1_EQ_1);
     if (B == 1'b0 && NCI1 == 1'b0)
       (A *> CO1) = (tpllh$A$CO1$B_EQ_0_AN_NCI1_EQ_0, tphhl$A$CO1$B_EQ_0_AN_NCI1_EQ_0);
     ifnone
       (A *> CO1) = (tpllh$A$CO1,tphhl$A$CO1);*/

// path delays
      (posedge A => (S +: S)) = (1.0, 1.0);
      (negedge A => (S -: S)) = (1.0, 1.0);
      if (B == 1'b1 && NCI1 == 1'b1) (A +=> CO1) = (1.0, 1.0);
      if (B == 1'b0 && NCI1 == 1'b0) (A +=> CO1) = (1.0, 1.0);

      if (B == 1'b1 && NCI2 == 1'b0) (A +=> CO2) = (1.0, 1.0);
      if (B == 1'b0 && NCI2 == 1'b0) (A +=> CO2) = (1.0, 1.0);


      if (B == 1'b1 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b0) (A +=> S) = (1.0, 1.0);
      if (B == 1'b1 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b1) (A +=> S) = (1.0, 1.0);
      if (B == 1'b1 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b0) (A +=> S) = (1.0, 1.0);
      if (B == 1'b0 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b1) (A +=> S) = (1.0, 1.0);
      if (B == 1'b0 && CS == 1'b1 && NCI1 == 1'b0 && NCI2 == 1'b1) (A +=> S) = (1.0, 1.0);
      if (B == 1'b0 && CS == 1'b0 && NCI1 == 1'b1 && NCI2 == 1'b0) (A +=> S) = (1.0, 1.0);
   

      if (B == 1'b0 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b0) (A -=> S) = (1.0, 1.0);
      if (B == 1'b0 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b1) (A -=> S) = (1.0, 1.0);
      if (B == 1'b1 && CS == 1'b1 && NCI1 == 1'b0 && NCI2 == 1'b1) (A -=> S) = (1.0, 1.0);
      if (B == 1'b1 && CS == 1'b0 && NCI1 == 1'b1 && NCI2 == 1'b0) (A -=> S) = (1.0, 1.0);
      if (B == 1'b1 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b1) (A -=> S) = (1.0, 1.0);
      if (B == 1'b0 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b0) (A -=> S) = (1.0, 1.0);

      (posedge B => (S +: S)) = (1.0, 1.0);
      (negedge B => (S -: S)) = (1.0, 1.0);
      if (A == 1'b1 && NCI1 == 1'b1) (B +=> CO1) = (1.0, 1.0);
      if (A == 1'b0 && NCI1 == 1'b0) (B +=> CO1) = (1.0, 1.0);
  
      if (A == 1'b1 && NCI2 == 1'b1) (B +=> CO2) = (1.0, 1.0);
      if (A == 1'b0 && NCI2 == 1'b0) (B +=> CO2) = (1.0, 1.0);
  

      if (A == 1'b1 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b0) (B +=> S) = (1.0, 1.0);
      if (A == 1'b1 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b1) (B +=> S) = (1.0, 1.0);
      if (A == 1'b1 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b0) (B +=> S) = (1.0, 1.0);
      if (A == 1'b0 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b1) (B +=> S) = (1.0, 1.0);
      if (A == 1'b0 && CS == 1'b1 && NCI1 == 1'b0 && NCI2 == 1'b1) (B +=> S) = (1.0, 1.0);
      if (A == 1'b0 && CS == 1'b0 && NCI1 == 1'b1 && NCI2 == 1'b0) (B +=> S) = (1.0, 1.0);
   

      if (A == 1'b0 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b0) (B -=> S) = (1.0, 1.0);
      if (A == 1'b0 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b1) (B -=> S) = (1.0, 1.0);
      if (A == 1'b1 && CS == 1'b1 && NCI1 == 1'b0 && NCI2 == 1'b1) (B -=> S) = (1.0, 1.0);
      if (A == 1'b1 && CS == 1'b0 && NCI1 == 1'b1 && NCI2 == 1'b0) (B -=> S) = (1.0, 1.0);
      if (A == 1'b1 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b1) (B -=> S) = (1.0, 1.0);
      if (A == 1'b0 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b0) (B -=> S) = (1.0, 1.0);


      (posedge NCI1 => (S +: S)) = (1.0, 1.0);
      (negedge NCI1 => (S -: S)) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1) (NCI1 -=> CO1) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0) (NCI1 -=> CO1) = (1.0, 1.0);

      
      if (A == 1'b1 && B == 1'b0 && CS == 1'b0 && NCI2 == 1'b1) (NCI1 +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1 && CS == 1'b0 && NCI2 == 1'b1) (NCI1 +=> S) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0 && CS == 1'b0 && NCI2 == 1'b0) (NCI1 +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1 && CS == 1'b0 && NCI2 == 1'b0) (NCI1 +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b0 && CS == 1'b0 && NCI2 == 1'b0) (NCI1 -=> S) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b1 && CS == 1'b0 && NCI2 == 1'b1) (NCI1 -=> S) = (1.0, 1.0);
   

      (posedge NCI2 => (S +: S)) = (1.0, 1.0);
      (negedge NCI2 => (S -: S)) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1) (NCI2 -=> CO2) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0) (NCI2 -=> CO2) = (1.0, 1.0);

      if (A == 1'b1 && B == 1'b0 && CS == 1'b1 && NCI1 == 1'b1) (NCI2 +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1 && CS == 1'b1 && NCI1 == 1'b1) (NCI2 +=> S) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0 && CS == 1'b1 && NCI1 == 1'b0) (NCI2 +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1 && CS == 1'b1 && NCI1 == 1'b0) (NCI2 +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b0 && CS == 1'b1 && NCI1 == 1'b0) (NCI2 -=> S) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b1 && CS == 1'b1 && NCI1 == 1'b1) (NCI2 -=> S) = (1.0, 1.0);

      (posedge CS => (S +: S)) = (1.0, 1.0);
      (negedge CS => (S -: S)) = (1.0, 1.0);

      if (A == 1'b1 && B == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b0) (CS +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b0 && NCI1 == 1'b1 && NCI2 == 1'b0) (CS +=> S) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b1 && NCI1 == 1'b0 && NCI2 == 1'b1) (CS -=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b1) (CS -=> S) = (1.0, 1.0);


   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_FA05D2 (CO1, CO2, S, A, B, CS, NCI1, NCI2);
input  A ;
input  B ;
input  CS ;
input  NCI1 ;
input  NCI2 ;
output CO1 ;
output CO2 ;
output S ;

   not (I0_out, NCI1);
   and (I1_out, I0_out, A);
   and (I2_out, A, B);
   not (I4_out, NCI1);
   and (I5_out, B, I4_out);
   or  (CO1, I1_out, I2_out, I5_out);
   not (I7_out, NCI2);
   and (I8_out, I7_out, A);
   and (I9_out, A, B);
   not (I11_out, NCI2);
   and (I12_out, B, I11_out);
   or  (CO2, I8_out, I9_out, I12_out);
   udp_mux2 (I14_out, NCI1, NCI2, CS);
   xor (I15_out, I14_out, A);
   xor (I16_out, I15_out, B);
   not (S, I16_out);

   specify
     // delay parameters
  /*   specparam
       tpllh$A$CO1 = 1.0,
       tphhl$A$CO1 = 1.0,
       tpllh$A$CO2 = 1.0,
       tphhl$A$CO2 = 1.0,
       tpllh$A$S = 1.0,
       tplhl$A$S = 1.0,
       tphlh$A$S = 1.0,
       tphhl$A$S = 1.0,
       tpllh$B$CO1 = 1.0,
       tphhl$B$CO1 = 1.0,
       tpllh$B$CO2 = 1.0,
       tphhl$B$CO2 = 1.0,
       tpllh$B$S = 1.0,
       tplhl$B$S = 1.0,
       tphlh$B$S = 1.0,
       tphhl$B$S = 1.0,
       tpllh$CS$S = 1.0,
       tplhl$CS$S = 1.0,
       tphlh$CS$S = 1.0,
       tphhl$CS$S = 1.0,
       tpllh$NCI1$S = 1.0,
       tplhl$NCI1$S = 1.0,
       tphlh$NCI1$S = 1.0,
       tphhl$NCI1$S = 1.0,
       tplhl$NCI1$CO1 = 1.0,
       tphlh$NCI1$CO1 = 1.0,
       tpllh$NCI2$S = 1.0,
       tplhl$NCI2$S = 1.0,
       tphlh$NCI2$S = 1.0,
       tphhl$NCI2$S = 1.0,
       tplhl$NCI2$CO2 = 1.0,
       tphlh$NCI2$CO2 = 1.0,
       tpllh$A$CO1$B_EQ_1_AN_NCI1_EQ_1 = 1.0,
       tphhl$A$CO1$B_EQ_1_AN_NCI1_EQ_1 = 1.0,
       tpllh$A$CO1$B_EQ_0_AN_NCI1_EQ_0 = 1.0,
       tphhl$A$CO1$B_EQ_0_AN_NCI1_EQ_0 = 1.0,
       tpllh$A$CO2$B_EQ_1_AN_NCI2_EQ_1 = 1.0,
       tphhl$A$CO2$B_EQ_1_AN_NCI2_EQ_1 = 1.0,
       tpllh$A$CO2$B_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tphhl$A$CO2$B_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tpllh$A$S$B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tphhl$A$S$B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tpllh$A$S$B_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tphhl$A$S$B_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tpllh$A$S$B_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tphhl$A$S$B_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tpllh$A$S$B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1 = 1.0,
       tphhl$A$S$B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1 = 1.0,
       tpllh$A$S$B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tphhl$A$S$B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tpllh$A$S$B_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tphhl$A$S$B_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tplhl$A$S$B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tphlh$A$S$B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tplhl$A$S$B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tphlh$A$S$B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tplhl$A$S$B_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tphlh$A$S$B_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tplhl$A$S$B_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tphlh$A$S$B_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tplhl$A$S$B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1 = 1.0,
       tphlh$A$S$B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1 = 1.0,
       tplhl$A$S$B_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tphlh$A$S$B_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tpllh$B$CO1$A_EQ_1_AN_NCI1_EQ_1 = 1.0,
       tphhl$B$CO1$A_EQ_1_AN_NCI1_EQ_1 = 1.0,
       tpllh$B$CO1$A_EQ_0_AN_NCI1_EQ_0 = 1.0,
       tphhl$B$CO1$A_EQ_0_AN_NCI1_EQ_0 = 1.0,
       tpllh$B$CO2$A_EQ_1_AN_NCI2_EQ_1 = 1.0,
       tphhl$B$CO2$A_EQ_1_AN_NCI2_EQ_1 = 1.0,
       tpllh$B$CO2$A_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tphhl$B$CO2$A_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tpllh$B$S$A_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tphhl$B$S$A_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tpllh$B$S$A_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tphhl$B$S$A_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tpllh$B$S$A_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tphhl$B$S$A_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tpllh$B$S$A_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1 = 1.0,
       tphhl$B$S$A_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1 = 1.0,
       tpllh$B$S$A_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tphhl$B$S$A_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tpllh$B$S$A_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tphhl$B$S$A_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tplhl$B$S$A_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tphlh$B$S$A_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tplhl$B$S$A_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tphlh$B$S$A_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tplhl$B$S$A_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tphlh$B$S$A_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tplhl$B$S$A_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tphlh$B$S$A_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tplhl$B$S$A_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1 = 1.0,
       tphlh$B$S$A_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1 = 1.0,
       tplhl$B$S$A_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tphlh$B$S$A_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tpllh$CS$S$A_EQ_1_AN_B_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tphhl$CS$S$A_EQ_1_AN_B_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tpllh$CS$S$A_EQ_0_AN_B_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tphhl$CS$S$A_EQ_0_AN_B_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tplhl$CS$S$A_EQ_0_AN_B_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tphlh$CS$S$A_EQ_0_AN_B_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tplhl$CS$S$A_EQ_1_AN_B_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tphlh$CS$S$A_EQ_1_AN_B_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tpllh$NCI1$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tphhl$NCI1$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tpllh$NCI1$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tphhl$NCI1$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tpllh$NCI1$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tphhl$NCI1$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tpllh$NCI1$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tphhl$NCI1$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tplhl$NCI1$S$A_EQ_0_AN_B_EQ_0_AN_CS_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tphlh$NCI1$S$A_EQ_0_AN_B_EQ_0_AN_CS_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tplhl$NCI1$S$A_EQ_1_AN_B_EQ_1_AN_CS_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tphlh$NCI1$S$A_EQ_1_AN_B_EQ_1_AN_CS_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tplhl$NCI1$CO1$A_EQ_0_AN_B_EQ_1 = 1.0,
       tphlh$NCI1$CO1$A_EQ_0_AN_B_EQ_1 = 1.0,
       tplhl$NCI1$CO1$A_EQ_1_AN_B_EQ_0 = 1.0,
       tphlh$NCI1$CO1$A_EQ_1_AN_B_EQ_0 = 1.0,
       tpllh$NCI2$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1 = 1.0,
       tphhl$NCI2$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1 = 1.0,
       tpllh$NCI2$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1 = 1.0,
       tphhl$NCI2$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1 = 1.0,
       tpllh$NCI2$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0 = 1.0,
       tphhl$NCI2$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0 = 1.0,
       tpllh$NCI2$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_0 = 1.0,
       tphhl$NCI2$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_0 = 1.0,
       tplhl$NCI2$S$A_EQ_0_AN_B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0 = 1.0,
       tphlh$NCI2$S$A_EQ_0_AN_B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0 = 1.0,
       tplhl$NCI2$S$A_EQ_1_AN_B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1 = 1.0,
       tphlh$NCI2$S$A_EQ_1_AN_B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1 = 1.0,
       tplhl$NCI2$CO2$A_EQ_0_AN_B_EQ_1 = 1.0,
       tphlh$NCI2$CO2$A_EQ_0_AN_B_EQ_1 = 1.0,
       tplhl$NCI2$CO2$A_EQ_1_AN_B_EQ_0 = 1.0,
       tphlh$NCI2$CO2$A_EQ_1_AN_B_EQ_0 = 1.0;

     // path delays
     if (A == 1'b1 && B == 1'b1 && CS == 1'b1 && NCI1 == 1'b1)
       (NCI2 *> S) = (tphlh$NCI2$S$A_EQ_1_AN_B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1, tplhl$NCI2$S$A_EQ_1_AN_B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1);
     if (A == 1'b1 && B == 1'b0 && CS == 1'b1 && NCI1 == 1'b1)
       (NCI2 *> S) = (tpllh$NCI2$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1, tphhl$NCI2$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1);
     if (A == 1'b1 && B == 1'b0 && CS == 1'b1 && NCI1 == 1'b0)
       (NCI2 *> S) = (tpllh$NCI2$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0, tphhl$NCI2$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0);
     if (A == 1'b0 && B == 1'b1 && CS == 1'b1 && NCI1 == 1'b1)
       (NCI2 *> S) = (tpllh$NCI2$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1, tphhl$NCI2$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1);
     if (A == 1'b0 && B == 1'b1 && CS == 1'b1 && NCI1 == 1'b0)
       (NCI2 *> S) = (tpllh$NCI2$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_0, tphhl$NCI2$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_0);
     if (A == 1'b0 && B == 1'b0 && CS == 1'b1 && NCI1 == 1'b0)
       (NCI2 *> S) = (tphlh$NCI2$S$A_EQ_0_AN_B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0, tplhl$NCI2$S$A_EQ_0_AN_B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0);
     ifnone
       (NCI2 *> S) = (tpllh$NCI2$S,tplhl$NCI2$S);

     if (A == 1'b1 && B == 1'b0)
       (NCI2 *> CO2) = (tphlh$NCI2$CO2$A_EQ_1_AN_B_EQ_0, tplhl$NCI2$CO2$A_EQ_1_AN_B_EQ_0);
     if (A == 1'b0 && B == 1'b1)
       (NCI2 *> CO2) = (tphlh$NCI2$CO2$A_EQ_0_AN_B_EQ_1, tplhl$NCI2$CO2$A_EQ_0_AN_B_EQ_1);
     ifnone
       (NCI2 *> CO2) = (tphlh$NCI2$CO2,tplhl$NCI2$CO2);

     if (A == 1'b1 && B == 1'b1 && CS == 1'b0 && NCI2 == 1'b1)
       (NCI1 *> S) = (tphlh$NCI1$S$A_EQ_1_AN_B_EQ_1_AN_CS_EQ_0_AN_NCI2_EQ_1, tplhl$NCI1$S$A_EQ_1_AN_B_EQ_1_AN_CS_EQ_0_AN_NCI2_EQ_1);
     if (A == 1'b1 && B == 1'b0 && CS == 1'b0 && NCI2 == 1'b1)
       (NCI1 *> S) = (tpllh$NCI1$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_0_AN_NCI2_EQ_1, tphhl$NCI1$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_0_AN_NCI2_EQ_1);
     if (A == 1'b1 && B == 1'b0 && CS == 1'b0 && NCI2 == 1'b0)
       (NCI1 *> S) = (tpllh$NCI1$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_0_AN_NCI2_EQ_0, tphhl$NCI1$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_0_AN_NCI2_EQ_0);
     if (A == 1'b0 && B == 1'b1 && CS == 1'b0 && NCI2 == 1'b1)
       (NCI1 *> S) = (tpllh$NCI1$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_0_AN_NCI2_EQ_1, tphhl$NCI1$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_0_AN_NCI2_EQ_1);
     if (A == 1'b0 && B == 1'b1 && CS == 1'b0 && NCI2 == 1'b0)
       (NCI1 *> S) = (tpllh$NCI1$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_0_AN_NCI2_EQ_0, tphhl$NCI1$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_0_AN_NCI2_EQ_0);
     if (A == 1'b0 && B == 1'b0 && CS == 1'b0 && NCI2 == 1'b0)
       (NCI1 *> S) = (tphlh$NCI1$S$A_EQ_0_AN_B_EQ_0_AN_CS_EQ_0_AN_NCI2_EQ_0, tplhl$NCI1$S$A_EQ_0_AN_B_EQ_0_AN_CS_EQ_0_AN_NCI2_EQ_0);
     ifnone
       (NCI1 *> S) = (tpllh$NCI1$S,tplhl$NCI1$S);

     if (A == 1'b1 && B == 1'b0)
       (NCI1 *> CO1) = (tphlh$NCI1$CO1$A_EQ_1_AN_B_EQ_0, tplhl$NCI1$CO1$A_EQ_1_AN_B_EQ_0);
     if (A == 1'b0 && B == 1'b1)
       (NCI1 *> CO1) = (tphlh$NCI1$CO1$A_EQ_0_AN_B_EQ_1, tplhl$NCI1$CO1$A_EQ_0_AN_B_EQ_1);
     ifnone
       (NCI1 *> CO1) = (tphlh$NCI1$CO1,tplhl$NCI1$CO1);

     if (A == 1'b1 && B == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b0)
       (CS *> S) = (tpllh$CS$S$A_EQ_1_AN_B_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0, tphhl$CS$S$A_EQ_1_AN_B_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0);
     if (A == 1'b1 && B == 1'b1 && NCI1 == 1'b0 && NCI2 == 1'b1)
       (CS *> S) = (tphlh$CS$S$A_EQ_1_AN_B_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1, tplhl$CS$S$A_EQ_1_AN_B_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1);
     if (A == 1'b0 && B == 1'b0 && NCI1 == 1'b1 && NCI2 == 1'b0)
       (CS *> S) = (tpllh$CS$S$A_EQ_0_AN_B_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0, tphhl$CS$S$A_EQ_0_AN_B_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0);
     if (A == 1'b0 && B == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b1)
       (CS *> S) = (tphlh$CS$S$A_EQ_0_AN_B_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1, tplhl$CS$S$A_EQ_0_AN_B_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1);
     ifnone
       (CS *> S) = (tpllh$CS$S,tplhl$CS$S);

     if (A == 1'b1 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b1)
       (B *> S) = (tphlh$B$S$A_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1, tplhl$B$S$A_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1);
     if (A == 1'b1 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b0)
       (B *> S) = (tpllh$B$S$A_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0, tphhl$B$S$A_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0);
     if (A == 1'b1 && CS == 1'b1 && NCI1 == 1'b0 && NCI2 == 1'b1)
       (B *> S) = (tphlh$B$S$A_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1, tplhl$B$S$A_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1);
     if (A == 1'b1 && CS == 1'b0 && NCI1 == 1'b1 && NCI2 == 1'b0)
       (B *> S) = (tphlh$B$S$A_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0, tplhl$B$S$A_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0);
     if (A == 1'b1 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b1)
       (B *> S) = (tpllh$B$S$A_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1, tphhl$B$S$A_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1);
     if (A == 1'b1 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b0)
       (B *> S) = (tpllh$B$S$A_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0, tphhl$B$S$A_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0);
     if (A == 1'b0 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b1)
       (B *> S) = (tpllh$B$S$A_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1, tphhl$B$S$A_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1);
     if (A == 1'b0 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b0)
       (B *> S) = (tphlh$B$S$A_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0, tplhl$B$S$A_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0);
     if (A == 1'b0 && CS == 1'b1 && NCI1 == 1'b0 && NCI2 == 1'b1)
       (B *> S) = (tpllh$B$S$A_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1, tphhl$B$S$A_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1);
     if (A == 1'b0 && CS == 1'b0 && NCI1 == 1'b1 && NCI2 == 1'b0)
       (B *> S) = (tpllh$B$S$A_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0, tphhl$B$S$A_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0);
     if (A == 1'b0 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b1)
       (B *> S) = (tphlh$B$S$A_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1, tplhl$B$S$A_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1);
     if (A == 1'b0 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b0)
       (B *> S) = (tphlh$B$S$A_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0, tplhl$B$S$A_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0);
     ifnone
       (B *> S) = (tpllh$B$S,tplhl$B$S);

     if (A == 1'b1 && NCI2 == 1'b1)
       (B *> CO2) = (tpllh$B$CO2$A_EQ_1_AN_NCI2_EQ_1, tphhl$B$CO2$A_EQ_1_AN_NCI2_EQ_1);
     if (A == 1'b0 && NCI2 == 1'b0)
       (B *> CO2) = (tpllh$B$CO2$A_EQ_0_AN_NCI2_EQ_0, tphhl$B$CO2$A_EQ_0_AN_NCI2_EQ_0);
     ifnone
       (B *> CO2) = (tpllh$B$CO2,tphhl$B$CO2);

     if (A == 1'b1 && NCI1 == 1'b1)
       (B *> CO1) = (tpllh$B$CO1$A_EQ_1_AN_NCI1_EQ_1, tphhl$B$CO1$A_EQ_1_AN_NCI1_EQ_1);
     if (A == 1'b0 && NCI1 == 1'b0)
       (B *> CO1) = (tpllh$B$CO1$A_EQ_0_AN_NCI1_EQ_0, tphhl$B$CO1$A_EQ_0_AN_NCI1_EQ_0);
     ifnone
       (B *> CO1) = (tpllh$B$CO1,tphhl$B$CO1);

     if (B == 1'b1 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b1)
       (A *> S) = (tphlh$A$S$B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1, tplhl$A$S$B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1);
     if (B == 1'b1 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b0)
       (A *> S) = (tpllh$A$S$B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0, tphhl$A$S$B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0);
     if (B == 1'b1 && CS == 1'b1 && NCI1 == 1'b0 && NCI2 == 1'b1)
       (A *> S) = (tphlh$A$S$B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1, tplhl$A$S$B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1);
     if (B == 1'b1 && CS == 1'b0 && NCI1 == 1'b1 && NCI2 == 1'b0)
       (A *> S) = (tphlh$A$S$B_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0, tplhl$A$S$B_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0);
     if (B == 1'b1 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b1)
       (A *> S) = (tpllh$A$S$B_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1, tphhl$A$S$B_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1);
     if (B == 1'b1 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b0)
       (A *> S) = (tpllh$A$S$B_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0, tphhl$A$S$B_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0);
     if (B == 1'b0 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b1)
       (A *> S) = (tpllh$A$S$B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1, tphhl$A$S$B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1);
     if (B == 1'b0 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b0)
       (A *> S) = (tphlh$A$S$B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0, tplhl$A$S$B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0);
     if (B == 1'b0 && CS == 1'b1 && NCI1 == 1'b0 && NCI2 == 1'b1)
       (A *> S) = (tpllh$A$S$B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1, tphhl$A$S$B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1);
     if (B == 1'b0 && CS == 1'b0 && NCI1 == 1'b1 && NCI2 == 1'b0)
       (A *> S) = (tpllh$A$S$B_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0, tphhl$A$S$B_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0);
     if (B == 1'b0 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b1)
       (A *> S) = (tphlh$A$S$B_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1, tplhl$A$S$B_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1);
     if (B == 1'b0 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b0)
       (A *> S) = (tphlh$A$S$B_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0, tplhl$A$S$B_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0);
     ifnone
       (A *> S) = (tpllh$A$S,tplhl$A$S);

     if (B == 1'b1 && NCI2 == 1'b1)
       (A *> CO2) = (tpllh$A$CO2$B_EQ_1_AN_NCI2_EQ_1, tphhl$A$CO2$B_EQ_1_AN_NCI2_EQ_1);
     if (B == 1'b0 && NCI2 == 1'b0)
       (A *> CO2) = (tpllh$A$CO2$B_EQ_0_AN_NCI2_EQ_0, tphhl$A$CO2$B_EQ_0_AN_NCI2_EQ_0);
     ifnone
       (A *> CO2) = (tpllh$A$CO2,tphhl$A$CO2);

     if (B == 1'b1 && NCI1 == 1'b1)
       (A *> CO1) = (tpllh$A$CO1$B_EQ_1_AN_NCI1_EQ_1, tphhl$A$CO1$B_EQ_1_AN_NCI1_EQ_1);
     if (B == 1'b0 && NCI1 == 1'b0)
       (A *> CO1) = (tpllh$A$CO1$B_EQ_0_AN_NCI1_EQ_0, tphhl$A$CO1$B_EQ_0_AN_NCI1_EQ_0);
     ifnone
       (A *> CO1) = (tpllh$A$CO1,tphhl$A$CO1);*/

// path delays
      (posedge A => (S +: S)) = (1.0, 1.0);
      (negedge A => (S -: S)) = (1.0, 1.0);
      if (B == 1'b1 && NCI1 == 1'b1) (A +=> CO1) = (1.0, 1.0);
      if (B == 1'b0 && NCI1 == 1'b0) (A +=> CO1) = (1.0, 1.0);

      if (B == 1'b1 && NCI2 == 1'b0) (A +=> CO2) = (1.0, 1.0);
      if (B == 1'b0 && NCI2 == 1'b0) (A +=> CO2) = (1.0, 1.0);


      if (B == 1'b1 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b0) (A +=> S) = (1.0, 1.0);
      if (B == 1'b1 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b1) (A +=> S) = (1.0, 1.0);
      if (B == 1'b1 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b0) (A +=> S) = (1.0, 1.0);
      if (B == 1'b0 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b1) (A +=> S) = (1.0, 1.0);
      if (B == 1'b0 && CS == 1'b1 && NCI1 == 1'b0 && NCI2 == 1'b1) (A +=> S) = (1.0, 1.0);
      if (B == 1'b0 && CS == 1'b0 && NCI1 == 1'b1 && NCI2 == 1'b0) (A +=> S) = (1.0, 1.0);
   

      if (B == 1'b0 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b0) (A -=> S) = (1.0, 1.0);
      if (B == 1'b0 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b1) (A -=> S) = (1.0, 1.0);
      if (B == 1'b1 && CS == 1'b1 && NCI1 == 1'b0 && NCI2 == 1'b1) (A -=> S) = (1.0, 1.0);
      if (B == 1'b1 && CS == 1'b0 && NCI1 == 1'b1 && NCI2 == 1'b0) (A -=> S) = (1.0, 1.0);
      if (B == 1'b1 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b1) (A -=> S) = (1.0, 1.0);
      if (B == 1'b0 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b0) (A -=> S) = (1.0, 1.0);

      (posedge B => (S +: S)) = (1.0, 1.0);
      (negedge B => (S -: S)) = (1.0, 1.0);
      if (A == 1'b1 && NCI1 == 1'b1) (B +=> CO1) = (1.0, 1.0);
      if (A == 1'b0 && NCI1 == 1'b0) (B +=> CO1) = (1.0, 1.0);
  
      if (A == 1'b1 && NCI2 == 1'b1) (B +=> CO2) = (1.0, 1.0);
      if (A == 1'b0 && NCI2 == 1'b0) (B +=> CO2) = (1.0, 1.0);
  

      if (A == 1'b1 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b0) (B +=> S) = (1.0, 1.0);
      if (A == 1'b1 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b1) (B +=> S) = (1.0, 1.0);
      if (A == 1'b1 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b0) (B +=> S) = (1.0, 1.0);
      if (A == 1'b0 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b1) (B +=> S) = (1.0, 1.0);
      if (A == 1'b0 && CS == 1'b1 && NCI1 == 1'b0 && NCI2 == 1'b1) (B +=> S) = (1.0, 1.0);
      if (A == 1'b0 && CS == 1'b0 && NCI1 == 1'b1 && NCI2 == 1'b0) (B +=> S) = (1.0, 1.0);
   

      if (A == 1'b0 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b0) (B -=> S) = (1.0, 1.0);
      if (A == 1'b0 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b1) (B -=> S) = (1.0, 1.0);
      if (A == 1'b1 && CS == 1'b1 && NCI1 == 1'b0 && NCI2 == 1'b1) (B -=> S) = (1.0, 1.0);
      if (A == 1'b1 && CS == 1'b0 && NCI1 == 1'b1 && NCI2 == 1'b0) (B -=> S) = (1.0, 1.0);
      if (A == 1'b1 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b1) (B -=> S) = (1.0, 1.0);
      if (A == 1'b0 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b0) (B -=> S) = (1.0, 1.0);


      (posedge NCI1 => (S +: S)) = (1.0, 1.0);
      (negedge NCI1 => (S -: S)) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1) (NCI1 -=> CO1) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0) (NCI1 -=> CO1) = (1.0, 1.0);

      
      if (A == 1'b1 && B == 1'b0 && CS == 1'b0 && NCI2 == 1'b1) (NCI1 +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1 && CS == 1'b0 && NCI2 == 1'b1) (NCI1 +=> S) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0 && CS == 1'b0 && NCI2 == 1'b0) (NCI1 +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1 && CS == 1'b0 && NCI2 == 1'b0) (NCI1 +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b0 && CS == 1'b0 && NCI2 == 1'b0) (NCI1 -=> S) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b1 && CS == 1'b0 && NCI2 == 1'b1) (NCI1 -=> S) = (1.0, 1.0);
   

      (posedge NCI2 => (S +: S)) = (1.0, 1.0);
      (negedge NCI2 => (S -: S)) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1) (NCI2 -=> CO2) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0) (NCI2 -=> CO2) = (1.0, 1.0);

      if (A == 1'b1 && B == 1'b0 && CS == 1'b1 && NCI1 == 1'b1) (NCI2 +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1 && CS == 1'b1 && NCI1 == 1'b1) (NCI2 +=> S) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0 && CS == 1'b1 && NCI1 == 1'b0) (NCI2 +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1 && CS == 1'b1 && NCI1 == 1'b0) (NCI2 +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b0 && CS == 1'b1 && NCI1 == 1'b0) (NCI2 -=> S) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b1 && CS == 1'b1 && NCI1 == 1'b1) (NCI2 -=> S) = (1.0, 1.0);

      (posedge CS => (S +: S)) = (1.0, 1.0);
      (negedge CS => (S -: S)) = (1.0, 1.0);

      if (A == 1'b1 && B == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b0) (CS +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b0 && NCI1 == 1'b1 && NCI2 == 1'b0) (CS +=> S) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b1 && NCI1 == 1'b0 && NCI2 == 1'b1) (CS -=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b1) (CS -=> S) = (1.0, 1.0);


   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_FA05D4 (CO1, CO2, S, A, B, CS, NCI1, NCI2);
input  A ;
input  B ;
input  CS ;
input  NCI1 ;
input  NCI2 ;
output CO1 ;
output CO2 ;
output S ;

   not (I0_out, NCI1);
   and (I1_out, I0_out, A);
   and (I2_out, A, B);
   not (I4_out, NCI1);
   and (I5_out, B, I4_out);
   or  (CO1, I1_out, I2_out, I5_out);
   not (I7_out, NCI2);
   and (I8_out, I7_out, A);
   and (I9_out, A, B);
   not (I11_out, NCI2);
   and (I12_out, B, I11_out);
   or  (CO2, I8_out, I9_out, I12_out);
   udp_mux2 (I14_out, NCI1, NCI2, CS);
   xor (I15_out, I14_out, A);
   xor (I16_out, I15_out, B);
   not (S, I16_out);

   specify
     // delay parameters
/*     specparam
       tpllh$A$CO1 = 1.0,
       tphhl$A$CO1 = 1.0,
       tpllh$A$CO2 = 1.0,
       tphhl$A$CO2 = 1.0,
       tpllh$A$S = 1.0,
       tplhl$A$S = 1.0,
       tphlh$A$S = 1.0,
       tphhl$A$S = 1.0,
       tpllh$B$CO1 = 1.0,
       tphhl$B$CO1 = 1.0,
       tpllh$B$CO2 = 1.0,
       tphhl$B$CO2 = 1.0,
       tpllh$B$S = 1.0,
       tplhl$B$S = 1.0,
       tphlh$B$S = 1.0,
       tphhl$B$S = 1.0,
       tpllh$CS$S = 1.0,
       tplhl$CS$S = 1.0,
       tphlh$CS$S = 1.0,
       tphhl$CS$S = 1.0,
       tpllh$NCI1$S = 1.0,
       tplhl$NCI1$S = 1.0,
       tphlh$NCI1$S = 1.0,
       tphhl$NCI1$S = 1.0,
       tplhl$NCI1$CO1 = 1.0,
       tphlh$NCI1$CO1 = 1.0,
       tpllh$NCI2$S = 1.0,
       tplhl$NCI2$S = 1.0,
       tphlh$NCI2$S = 1.0,
       tphhl$NCI2$S = 1.0,
       tplhl$NCI2$CO2 = 1.0,
       tphlh$NCI2$CO2 = 1.0,
       tpllh$A$CO1$B_EQ_1_AN_NCI1_EQ_1 = 1.0,
       tphhl$A$CO1$B_EQ_1_AN_NCI1_EQ_1 = 1.0,
       tpllh$A$CO1$B_EQ_0_AN_NCI1_EQ_0 = 1.0,
       tphhl$A$CO1$B_EQ_0_AN_NCI1_EQ_0 = 1.0,
       tpllh$A$CO2$B_EQ_1_AN_NCI2_EQ_1 = 1.0,
       tphhl$A$CO2$B_EQ_1_AN_NCI2_EQ_1 = 1.0,
       tpllh$A$CO2$B_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tphhl$A$CO2$B_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tpllh$A$S$B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tphhl$A$S$B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tpllh$A$S$B_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tphhl$A$S$B_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tpllh$A$S$B_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tphhl$A$S$B_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tpllh$A$S$B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1 = 1.0,
       tphhl$A$S$B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1 = 1.0,
       tpllh$A$S$B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tphhl$A$S$B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tpllh$A$S$B_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tphhl$A$S$B_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tplhl$A$S$B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tphlh$A$S$B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tplhl$A$S$B_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tphlh$A$S$B_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tplhl$A$S$B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1 = 1.0,
       tphlh$A$S$B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1 = 1.0,
       tplhl$A$S$B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tphlh$A$S$B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tplhl$A$S$B_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tphlh$A$S$B_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tplhl$A$S$B_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tphlh$A$S$B_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tpllh$B$CO1$A_EQ_1_AN_NCI1_EQ_1 = 1.0,
       tphhl$B$CO1$A_EQ_1_AN_NCI1_EQ_1 = 1.0,
       tpllh$B$CO1$A_EQ_0_AN_NCI1_EQ_0 = 1.0,
       tphhl$B$CO1$A_EQ_0_AN_NCI1_EQ_0 = 1.0,
       tpllh$B$CO2$A_EQ_1_AN_NCI2_EQ_1 = 1.0,
       tphhl$B$CO2$A_EQ_1_AN_NCI2_EQ_1 = 1.0,
       tpllh$B$CO2$A_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tphhl$B$CO2$A_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tpllh$B$S$A_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tphhl$B$S$A_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tpllh$B$S$A_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tphhl$B$S$A_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tpllh$B$S$A_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tphhl$B$S$A_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tpllh$B$S$A_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1 = 1.0,
       tphhl$B$S$A_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1 = 1.0,
       tpllh$B$S$A_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tphhl$B$S$A_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tpllh$B$S$A_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tphhl$B$S$A_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tplhl$B$S$A_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tphlh$B$S$A_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tplhl$B$S$A_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tphlh$B$S$A_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tplhl$B$S$A_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tphlh$B$S$A_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tplhl$B$S$A_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tphlh$B$S$A_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tplhl$B$S$A_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1 = 1.0,
       tphlh$B$S$A_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1 = 1.0,
       tplhl$B$S$A_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tphlh$B$S$A_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tpllh$CS$S$A_EQ_1_AN_B_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tphhl$CS$S$A_EQ_1_AN_B_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tpllh$CS$S$A_EQ_0_AN_B_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tphhl$CS$S$A_EQ_0_AN_B_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0 = 1.0,
       tplhl$CS$S$A_EQ_1_AN_B_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tphlh$CS$S$A_EQ_1_AN_B_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tplhl$CS$S$A_EQ_0_AN_B_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tphlh$CS$S$A_EQ_0_AN_B_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tpllh$NCI1$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tphhl$NCI1$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tpllh$NCI1$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tphhl$NCI1$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tpllh$NCI1$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tphhl$NCI1$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tpllh$NCI1$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tphhl$NCI1$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tplhl$NCI1$S$A_EQ_0_AN_B_EQ_0_AN_CS_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tphlh$NCI1$S$A_EQ_0_AN_B_EQ_0_AN_CS_EQ_0_AN_NCI2_EQ_0 = 1.0,
       tplhl$NCI1$S$A_EQ_1_AN_B_EQ_1_AN_CS_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tphlh$NCI1$S$A_EQ_1_AN_B_EQ_1_AN_CS_EQ_0_AN_NCI2_EQ_1 = 1.0,
       tplhl$NCI1$CO1$A_EQ_0_AN_B_EQ_1 = 1.0,
       tphlh$NCI1$CO1$A_EQ_0_AN_B_EQ_1 = 1.0,
       tplhl$NCI1$CO1$A_EQ_1_AN_B_EQ_0 = 1.0,
       tphlh$NCI1$CO1$A_EQ_1_AN_B_EQ_0 = 1.0,
       tpllh$NCI2$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1 = 1.0,
       tphhl$NCI2$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1 = 1.0,
       tpllh$NCI2$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1 = 1.0,
       tphhl$NCI2$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1 = 1.0,
       tpllh$NCI2$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_0 = 1.0,
       tphhl$NCI2$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_0 = 1.0,
       tpllh$NCI2$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0 = 1.0,
       tphhl$NCI2$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0 = 1.0,
       tplhl$NCI2$S$A_EQ_0_AN_B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0 = 1.0,
       tphlh$NCI2$S$A_EQ_0_AN_B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0 = 1.0,
       tplhl$NCI2$S$A_EQ_1_AN_B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1 = 1.0,
       tphlh$NCI2$S$A_EQ_1_AN_B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1 = 1.0,
       tplhl$NCI2$CO2$A_EQ_0_AN_B_EQ_1 = 1.0,
       tphlh$NCI2$CO2$A_EQ_0_AN_B_EQ_1 = 1.0,
       tplhl$NCI2$CO2$A_EQ_1_AN_B_EQ_0 = 1.0,
       tphlh$NCI2$CO2$A_EQ_1_AN_B_EQ_0 = 1.0;

     // path delays
     if (A == 1'b1 && B == 1'b1 && CS == 1'b1 && NCI1 == 1'b1)
       (NCI2 *> S) = (tphlh$NCI2$S$A_EQ_1_AN_B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1, tplhl$NCI2$S$A_EQ_1_AN_B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1);
     if (A == 1'b1 && B == 1'b0 && CS == 1'b1 && NCI1 == 1'b1)
       (NCI2 *> S) = (tpllh$NCI2$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1, tphhl$NCI2$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1);
     if (A == 1'b1 && B == 1'b0 && CS == 1'b1 && NCI1 == 1'b0)
       (NCI2 *> S) = (tpllh$NCI2$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0, tphhl$NCI2$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0);
     if (A == 1'b0 && B == 1'b1 && CS == 1'b1 && NCI1 == 1'b1)
       (NCI2 *> S) = (tpllh$NCI2$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1, tphhl$NCI2$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1);
     if (A == 1'b0 && B == 1'b1 && CS == 1'b1 && NCI1 == 1'b0)
       (NCI2 *> S) = (tpllh$NCI2$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_0, tphhl$NCI2$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_0);
     if (A == 1'b0 && B == 1'b0 && CS == 1'b1 && NCI1 == 1'b0)
       (NCI2 *> S) = (tphlh$NCI2$S$A_EQ_0_AN_B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0, tplhl$NCI2$S$A_EQ_0_AN_B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0);
     ifnone
       (NCI2 *> S) = (tpllh$NCI2$S,tplhl$NCI2$S);

     if (A == 1'b1 && B == 1'b0)
       (NCI2 *> CO2) = (tphlh$NCI2$CO2$A_EQ_1_AN_B_EQ_0, tplhl$NCI2$CO2$A_EQ_1_AN_B_EQ_0);
     if (A == 1'b0 && B == 1'b1)
       (NCI2 *> CO2) = (tphlh$NCI2$CO2$A_EQ_0_AN_B_EQ_1, tplhl$NCI2$CO2$A_EQ_0_AN_B_EQ_1);
     ifnone
       (NCI2 *> CO2) = (tphlh$NCI2$CO2,tplhl$NCI2$CO2);

     if (A == 1'b1 && B == 1'b1 && CS == 1'b0 && NCI2 == 1'b1)
       (NCI1 *> S) = (tphlh$NCI1$S$A_EQ_1_AN_B_EQ_1_AN_CS_EQ_0_AN_NCI2_EQ_1, tplhl$NCI1$S$A_EQ_1_AN_B_EQ_1_AN_CS_EQ_0_AN_NCI2_EQ_1);
     if (A == 1'b1 && B == 1'b0 && CS == 1'b0 && NCI2 == 1'b1)
       (NCI1 *> S) = (tpllh$NCI1$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_0_AN_NCI2_EQ_1, tphhl$NCI1$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_0_AN_NCI2_EQ_1);
     if (A == 1'b1 && B == 1'b0 && CS == 1'b0 && NCI2 == 1'b0)
       (NCI1 *> S) = (tpllh$NCI1$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_0_AN_NCI2_EQ_0, tphhl$NCI1$S$A_EQ_1_AN_B_EQ_0_AN_CS_EQ_0_AN_NCI2_EQ_0);
     if (A == 1'b0 && B == 1'b1 && CS == 1'b0 && NCI2 == 1'b1)
       (NCI1 *> S) = (tpllh$NCI1$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_0_AN_NCI2_EQ_1, tphhl$NCI1$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_0_AN_NCI2_EQ_1);
     if (A == 1'b0 && B == 1'b1 && CS == 1'b0 && NCI2 == 1'b0)
       (NCI1 *> S) = (tpllh$NCI1$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_0_AN_NCI2_EQ_0, tphhl$NCI1$S$A_EQ_0_AN_B_EQ_1_AN_CS_EQ_0_AN_NCI2_EQ_0);
     if (A == 1'b0 && B == 1'b0 && CS == 1'b0 && NCI2 == 1'b0)
       (NCI1 *> S) = (tphlh$NCI1$S$A_EQ_0_AN_B_EQ_0_AN_CS_EQ_0_AN_NCI2_EQ_0, tplhl$NCI1$S$A_EQ_0_AN_B_EQ_0_AN_CS_EQ_0_AN_NCI2_EQ_0);
     ifnone
       (NCI1 *> S) = (tpllh$NCI1$S,tplhl$NCI1$S);

     if (A == 1'b1 && B == 1'b0)
       (NCI1 *> CO1) = (tphlh$NCI1$CO1$A_EQ_1_AN_B_EQ_0, tplhl$NCI1$CO1$A_EQ_1_AN_B_EQ_0);
     if (A == 1'b0 && B == 1'b1)
       (NCI1 *> CO1) = (tphlh$NCI1$CO1$A_EQ_0_AN_B_EQ_1, tplhl$NCI1$CO1$A_EQ_0_AN_B_EQ_1);
     ifnone
       (NCI1 *> CO1) = (tphlh$NCI1$CO1,tplhl$NCI1$CO1);

     if (A == 1'b1 && B == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b0)
       (CS *> S) = (tpllh$CS$S$A_EQ_1_AN_B_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0, tphhl$CS$S$A_EQ_1_AN_B_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0);
     if (A == 1'b1 && B == 1'b1 && NCI1 == 1'b0 && NCI2 == 1'b1)
       (CS *> S) = (tphlh$CS$S$A_EQ_1_AN_B_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1, tplhl$CS$S$A_EQ_1_AN_B_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1);
     if (A == 1'b0 && B == 1'b0 && NCI1 == 1'b1 && NCI2 == 1'b0)
       (CS *> S) = (tpllh$CS$S$A_EQ_0_AN_B_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0, tphhl$CS$S$A_EQ_0_AN_B_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0);
     if (A == 1'b0 && B == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b1)
       (CS *> S) = (tphlh$CS$S$A_EQ_0_AN_B_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1, tplhl$CS$S$A_EQ_0_AN_B_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1);
     ifnone
       (CS *> S) = (tpllh$CS$S,tplhl$CS$S);

     if (A == 1'b1 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b1)
       (B *> S) = (tphlh$B$S$A_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1, tplhl$B$S$A_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1);
     if (A == 1'b1 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b0)
       (B *> S) = (tpllh$B$S$A_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0, tphhl$B$S$A_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0);
     if (A == 1'b1 && CS == 1'b1 && NCI1 == 1'b0 && NCI2 == 1'b1)
       (B *> S) = (tphlh$B$S$A_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1, tplhl$B$S$A_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1);
     if (A == 1'b1 && CS == 1'b0 && NCI1 == 1'b1 && NCI2 == 1'b0)
       (B *> S) = (tphlh$B$S$A_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0, tplhl$B$S$A_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0);
     if (A == 1'b1 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b1)
       (B *> S) = (tpllh$B$S$A_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1, tphhl$B$S$A_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1);
     if (A == 1'b1 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b0)
       (B *> S) = (tpllh$B$S$A_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0, tphhl$B$S$A_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0);
     if (A == 1'b0 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b1)
       (B *> S) = (tpllh$B$S$A_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1, tphhl$B$S$A_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1);
     if (A == 1'b0 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b0)
       (B *> S) = (tphlh$B$S$A_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0, tplhl$B$S$A_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0);
     if (A == 1'b0 && CS == 1'b1 && NCI1 == 1'b0 && NCI2 == 1'b1)
       (B *> S) = (tpllh$B$S$A_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1, tphhl$B$S$A_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1);
     if (A == 1'b0 && CS == 1'b0 && NCI1 == 1'b1 && NCI2 == 1'b0)
       (B *> S) = (tpllh$B$S$A_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0, tphhl$B$S$A_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0);
     if (A == 1'b0 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b1)
       (B *> S) = (tphlh$B$S$A_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1, tplhl$B$S$A_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1);
     if (A == 1'b0 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b0)
       (B *> S) = (tphlh$B$S$A_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0, tplhl$B$S$A_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0);
     ifnone
       (B *> S) = (tpllh$B$S,tplhl$B$S);

     if (A == 1'b1 && NCI2 == 1'b1)
       (B *> CO2) = (tpllh$B$CO2$A_EQ_1_AN_NCI2_EQ_1, tphhl$B$CO2$A_EQ_1_AN_NCI2_EQ_1);
     if (A == 1'b0 && NCI2 == 1'b0)
       (B *> CO2) = (tpllh$B$CO2$A_EQ_0_AN_NCI2_EQ_0, tphhl$B$CO2$A_EQ_0_AN_NCI2_EQ_0);
     ifnone
       (B *> CO2) = (tpllh$B$CO2,tphhl$B$CO2);

     if (A == 1'b1 && NCI1 == 1'b1)
       (B *> CO1) = (tpllh$B$CO1$A_EQ_1_AN_NCI1_EQ_1, tphhl$B$CO1$A_EQ_1_AN_NCI1_EQ_1);
     if (A == 1'b0 && NCI1 == 1'b0)
       (B *> CO1) = (tpllh$B$CO1$A_EQ_0_AN_NCI1_EQ_0, tphhl$B$CO1$A_EQ_0_AN_NCI1_EQ_0);
     ifnone
       (B *> CO1) = (tpllh$B$CO1,tphhl$B$CO1);

     if (B == 1'b1 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b1)
       (A *> S) = (tphlh$A$S$B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1, tplhl$A$S$B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1);
     if (B == 1'b1 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b0)
       (A *> S) = (tpllh$A$S$B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0, tphhl$A$S$B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0);
     if (B == 1'b1 && CS == 1'b1 && NCI1 == 1'b0 && NCI2 == 1'b1)
       (A *> S) = (tphlh$A$S$B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1, tplhl$A$S$B_EQ_1_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1);
     if (B == 1'b1 && CS == 1'b0 && NCI1 == 1'b1 && NCI2 == 1'b0)
       (A *> S) = (tphlh$A$S$B_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0, tplhl$A$S$B_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0);
     if (B == 1'b1 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b1)
       (A *> S) = (tpllh$A$S$B_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1, tphhl$A$S$B_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1);
     if (B == 1'b1 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b0)
       (A *> S) = (tpllh$A$S$B_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0, tphhl$A$S$B_EQ_1_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0);
     if (B == 1'b0 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b1)
       (A *> S) = (tpllh$A$S$B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1, tphhl$A$S$B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_1);
     if (B == 1'b0 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b0)
       (A *> S) = (tphlh$A$S$B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0, tplhl$A$S$B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_1_AN_NCI2_EQ_0);
     if (B == 1'b0 && CS == 1'b1 && NCI1 == 1'b0 && NCI2 == 1'b1)
       (A *> S) = (tpllh$A$S$B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1, tphhl$A$S$B_EQ_0_AN_CS_EQ_1_AN_NCI1_EQ_0_AN_NCI2_EQ_1);
     if (B == 1'b0 && CS == 1'b0 && NCI1 == 1'b1 && NCI2 == 1'b0)
       (A *> S) = (tpllh$A$S$B_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0, tphhl$A$S$B_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_1_AN_NCI2_EQ_0);
     if (B == 1'b0 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b1)
       (A *> S) = (tphlh$A$S$B_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1, tplhl$A$S$B_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_1);
     if (B == 1'b0 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b0)
       (A *> S) = (tphlh$A$S$B_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0, tplhl$A$S$B_EQ_0_AN_CS_EQ_0_AN_NCI1_EQ_0_AN_NCI2_EQ_0);
     ifnone
       (A *> S) = (tpllh$A$S,tplhl$A$S);

     if (B == 1'b1 && NCI2 == 1'b1)
       (A *> CO2) = (tpllh$A$CO2$B_EQ_1_AN_NCI2_EQ_1, tphhl$A$CO2$B_EQ_1_AN_NCI2_EQ_1);
     if (B == 1'b0 && NCI2 == 1'b0)
       (A *> CO2) = (tpllh$A$CO2$B_EQ_0_AN_NCI2_EQ_0, tphhl$A$CO2$B_EQ_0_AN_NCI2_EQ_0);
     ifnone
       (A *> CO2) = (tpllh$A$CO2,tphhl$A$CO2);

     if (B == 1'b1 && NCI1 == 1'b1)
       (A *> CO1) = (tpllh$A$CO1$B_EQ_1_AN_NCI1_EQ_1, tphhl$A$CO1$B_EQ_1_AN_NCI1_EQ_1);
     if (B == 1'b0 && NCI1 == 1'b0)
       (A *> CO1) = (tpllh$A$CO1$B_EQ_0_AN_NCI1_EQ_0, tphhl$A$CO1$B_EQ_0_AN_NCI1_EQ_0);
     ifnone
       (A *> CO1) = (tpllh$A$CO1,tphhl$A$CO1);*/

// path delays
      (posedge A => (S +: S)) = (1.0, 1.0);
      (negedge A => (S -: S)) = (1.0, 1.0);
      if (B == 1'b1 && NCI1 == 1'b1) (A +=> CO1) = (1.0, 1.0);
      if (B == 1'b0 && NCI1 == 1'b0) (A +=> CO1) = (1.0, 1.0);

      if (B == 1'b1 && NCI2 == 1'b0) (A +=> CO2) = (1.0, 1.0);
      if (B == 1'b0 && NCI2 == 1'b0) (A +=> CO2) = (1.0, 1.0);


      if (B == 1'b1 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b0) (A +=> S) = (1.0, 1.0);
      if (B == 1'b1 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b1) (A +=> S) = (1.0, 1.0);
      if (B == 1'b1 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b0) (A +=> S) = (1.0, 1.0);
      if (B == 1'b0 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b1) (A +=> S) = (1.0, 1.0);
      if (B == 1'b0 && CS == 1'b1 && NCI1 == 1'b0 && NCI2 == 1'b1) (A +=> S) = (1.0, 1.0);
      if (B == 1'b0 && CS == 1'b0 && NCI1 == 1'b1 && NCI2 == 1'b0) (A +=> S) = (1.0, 1.0);
   

      if (B == 1'b0 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b0) (A -=> S) = (1.0, 1.0);
      if (B == 1'b0 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b1) (A -=> S) = (1.0, 1.0);
      if (B == 1'b1 && CS == 1'b1 && NCI1 == 1'b0 && NCI2 == 1'b1) (A -=> S) = (1.0, 1.0);
      if (B == 1'b1 && CS == 1'b0 && NCI1 == 1'b1 && NCI2 == 1'b0) (A -=> S) = (1.0, 1.0);
      if (B == 1'b1 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b1) (A -=> S) = (1.0, 1.0);
      if (B == 1'b0 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b0) (A -=> S) = (1.0, 1.0);

      (posedge B => (S +: S)) = (1.0, 1.0);
      (negedge B => (S -: S)) = (1.0, 1.0);
      if (A == 1'b1 && NCI1 == 1'b1) (B +=> CO1) = (1.0, 1.0);
      if (A == 1'b0 && NCI1 == 1'b0) (B +=> CO1) = (1.0, 1.0);
  
      if (A == 1'b1 && NCI2 == 1'b1) (B +=> CO2) = (1.0, 1.0);
      if (A == 1'b0 && NCI2 == 1'b0) (B +=> CO2) = (1.0, 1.0);
  

      if (A == 1'b1 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b0) (B +=> S) = (1.0, 1.0);
      if (A == 1'b1 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b1) (B +=> S) = (1.0, 1.0);
      if (A == 1'b1 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b0) (B +=> S) = (1.0, 1.0);
      if (A == 1'b0 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b1) (B +=> S) = (1.0, 1.0);
      if (A == 1'b0 && CS == 1'b1 && NCI1 == 1'b0 && NCI2 == 1'b1) (B +=> S) = (1.0, 1.0);
      if (A == 1'b0 && CS == 1'b0 && NCI1 == 1'b1 && NCI2 == 1'b0) (B +=> S) = (1.0, 1.0);
   

      if (A == 1'b0 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b0) (B -=> S) = (1.0, 1.0);
      if (A == 1'b0 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b1) (B -=> S) = (1.0, 1.0);
      if (A == 1'b1 && CS == 1'b1 && NCI1 == 1'b0 && NCI2 == 1'b1) (B -=> S) = (1.0, 1.0);
      if (A == 1'b1 && CS == 1'b0 && NCI1 == 1'b1 && NCI2 == 1'b0) (B -=> S) = (1.0, 1.0);
      if (A == 1'b1 && CS == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b1) (B -=> S) = (1.0, 1.0);
      if (A == 1'b0 && CS == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b0) (B -=> S) = (1.0, 1.0);


      (posedge NCI1 => (S +: S)) = (1.0, 1.0);
      (negedge NCI1 => (S -: S)) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1) (NCI1 -=> CO1) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0) (NCI1 -=> CO1) = (1.0, 1.0);

      
      if (A == 1'b1 && B == 1'b0 && CS == 1'b0 && NCI2 == 1'b1) (NCI1 +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1 && CS == 1'b0 && NCI2 == 1'b1) (NCI1 +=> S) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0 && CS == 1'b0 && NCI2 == 1'b0) (NCI1 +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1 && CS == 1'b0 && NCI2 == 1'b0) (NCI1 +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b0 && CS == 1'b0 && NCI2 == 1'b0) (NCI1 -=> S) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b1 && CS == 1'b0 && NCI2 == 1'b1) (NCI1 -=> S) = (1.0, 1.0);
   

      (posedge NCI2 => (S +: S)) = (1.0, 1.0);
      (negedge NCI2 => (S -: S)) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1) (NCI2 -=> CO2) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0) (NCI2 -=> CO2) = (1.0, 1.0);

      if (A == 1'b1 && B == 1'b0 && CS == 1'b1 && NCI1 == 1'b1) (NCI2 +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1 && CS == 1'b1 && NCI1 == 1'b1) (NCI2 +=> S) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b0 && CS == 1'b1 && NCI1 == 1'b0) (NCI2 +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b1 && CS == 1'b1 && NCI1 == 1'b0) (NCI2 +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b0 && CS == 1'b1 && NCI1 == 1'b0) (NCI2 -=> S) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b1 && CS == 1'b1 && NCI1 == 1'b1) (NCI2 -=> S) = (1.0, 1.0);

      (posedge CS => (S +: S)) = (1.0, 1.0);
      (negedge CS => (S -: S)) = (1.0, 1.0);

      if (A == 1'b1 && B == 1'b1 && NCI1 == 1'b1 && NCI2 == 1'b0) (CS +=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b0 && NCI1 == 1'b1 && NCI2 == 1'b0) (CS +=> S) = (1.0, 1.0);
      if (A == 1'b1 && B == 1'b1 && NCI1 == 1'b0 && NCI2 == 1'b1) (CS -=> S) = (1.0, 1.0);
      if (A == 1'b0 && B == 1'b0 && NCI1 == 1'b0 && NCI2 == 1'b1) (CS -=> S) = (1.0, 1.0);


   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_FVDD (Z);
output Z ;

   buf (Z, 1'B1);


endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_FVSS (Z);
output Z ;

   buf (Z, 1'B0);


endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_HA01D1 (CO, S, A, B);
input  A ;
input  B ;
output CO ;
output S ;

   and (CO, A, B);
   xor (S, A, B);

   specify
     // delay parameters
     specparam
       tpllh$A$S = 1.0,
       tplhl$A$S = 1.0,
       tphlh$A$S = 1.0,
       tphhl$A$S = 1.0,
       tpllh$A$CO = 1.0,
       tphhl$A$CO = 1.0,
       tpllh$B$S = 1.0,
       tplhl$B$S = 1.0,
       tphlh$B$S = 1.0,
       tphhl$B$S = 1.0,
       tpllh$B$CO = 1.0,
       tphhl$B$CO = 1.0;

     // path delays
     (posedge B *> (S +: !A)) = (tpllh$B$S, tplhl$B$S);
     (negedge B *> (S +: A)) = (tphlh$B$S, tphhl$B$S);
     (B *> CO) = (tpllh$B$CO, tphhl$B$CO);
     (posedge A *> (S +: !B)) = (tpllh$A$S, tplhl$A$S);
     (negedge A *> (S +: B)) = (tphlh$A$S, tphhl$A$S);
     (A *> CO) = (tpllh$A$CO, tphhl$A$CO);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_HA01D2 (CO, S, A, B);
input  A ;
input  B ;
output CO ;
output S ;

   and (CO, A, B);
   xor (S, A, B);

   specify
     // delay parameters
     specparam
       tpllh$A$S = 1.0,
       tplhl$A$S = 1.0,
       tphlh$A$S = 1.0,
       tphhl$A$S = 1.0,
       tpllh$A$CO = 1.0,
       tphhl$A$CO = 1.0,
       tpllh$B$S = 1.0,
       tplhl$B$S = 1.0,
       tphlh$B$S = 1.0,
       tphhl$B$S = 1.0,
       tpllh$B$CO = 1.0,
       tphhl$B$CO = 1.0;

     // path delays
     (posedge B *> (S +: !A)) = (tpllh$B$S, tplhl$B$S);
     (negedge B *> (S +: A)) = (tphlh$B$S, tphhl$B$S);
     (B *> CO) = (tpllh$B$CO, tphhl$B$CO);
     (posedge A *> (S +: !B)) = (tpllh$A$S, tplhl$A$S);
     (negedge A *> (S +: B)) = (tphlh$A$S, tphhl$A$S);
     (A *> CO) = (tpllh$A$CO, tphhl$A$CO);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_HA01D4 (CO, S, A, B);
input  A ;
input  B ;
output CO ;
output S ;

   and (CO, A, B);
   xor (S, A, B);

   specify
     // delay parameters
     specparam
       tpllh$A$S = 1.0,
       tplhl$A$S = 1.0,
       tphlh$A$S = 1.0,
       tphhl$A$S = 1.0,
       tpllh$A$CO = 1.0,
       tphhl$A$CO = 1.0,
       tpllh$B$S = 1.0,
       tplhl$B$S = 1.0,
       tphlh$B$S = 1.0,
       tphhl$B$S = 1.0,
       tpllh$B$CO = 1.0,
       tphhl$B$CO = 1.0;

     // path delays
     (posedge B *> (S +: !A)) = (tpllh$B$S, tplhl$B$S);
     (negedge B *> (S +: A)) = (tphlh$B$S, tphhl$B$S);
     (B *> CO) = (tpllh$B$CO, tphhl$B$CO);
     (posedge A *> (S +: !B)) = (tpllh$A$S, tplhl$A$S);
     (negedge A *> (S +: B)) = (tphlh$A$S, tphhl$A$S);
     (A *> CO) = (tpllh$A$CO, tphhl$A$CO);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_HA02D1 (NCO, S, A, CI);
input  A ;
input  CI ;
output NCO ;
output S ;

   and (I0_out, A, CI);
   not (NCO, I0_out);
   xor (S, A, CI);

   specify
     // delay parameters
     specparam
       tpllh$A$S = 1.0,
       tplhl$A$S = 1.0,
       tphlh$A$S = 1.0,
       tphhl$A$S = 1.0,
       tplhl$A$NCO = 1.0,
       tphlh$A$NCO = 1.0,
       tpllh$CI$S = 1.0,
       tplhl$CI$S = 1.0,
       tphlh$CI$S = 1.0,
       tphhl$CI$S = 1.0,
       tplhl$CI$NCO = 1.0,
       tphlh$CI$NCO = 1.0;

     // path delays
     (posedge CI *> (S +: !A)) = (tpllh$CI$S, tplhl$CI$S);
     (negedge CI *> (S +: A)) = (tphlh$CI$S, tphhl$CI$S);
     (CI *> NCO) = (tphlh$CI$NCO, tplhl$CI$NCO);
     (posedge A *> (S +: !CI)) = (tpllh$A$S, tplhl$A$S);
     (negedge A *> (S +: CI)) = (tphlh$A$S, tphhl$A$S);
     (A *> NCO) = (tphlh$A$NCO, tplhl$A$NCO);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_HA02D2 (NCO, S, A, CI);
input  A ;
input  CI ;
output NCO ;
output S ;

   and (I0_out, A, CI);
   not (NCO, I0_out);
   xor (S, A, CI);

   specify
     // delay parameters
     specparam
       tpllh$A$S = 1.0,
       tplhl$A$S = 1.0,
       tphlh$A$S = 1.0,
       tphhl$A$S = 1.0,
       tplhl$A$NCO = 1.0,
       tphlh$A$NCO = 1.0,
       tpllh$CI$S = 1.0,
       tplhl$CI$S = 1.0,
       tphlh$CI$S = 1.0,
       tphhl$CI$S = 1.0,
       tplhl$CI$NCO = 1.0,
       tphlh$CI$NCO = 1.0;

     // path delays
     (posedge CI *> (S +: !A)) = (tpllh$CI$S, tplhl$CI$S);
     (negedge CI *> (S +: A)) = (tphlh$CI$S, tphhl$CI$S);
     (CI *> NCO) = (tphlh$CI$NCO, tplhl$CI$NCO);
     (posedge A *> (S +: !CI)) = (tpllh$A$S, tplhl$A$S);
     (negedge A *> (S +: CI)) = (tphlh$A$S, tphhl$A$S);
     (A *> NCO) = (tphlh$A$NCO, tplhl$A$NCO);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_HA02D4 (NCO, S, A, CI);
input  A ;
input  CI ;
output NCO ;
output S ;

   and (I0_out, A, CI);
   not (NCO, I0_out);
   xor (S, A, CI);

   specify
     // delay parameters
     specparam
       tpllh$A$S = 1.0,
       tplhl$A$S = 1.0,
       tphlh$A$S = 1.0,
       tphhl$A$S = 1.0,
       tplhl$A$NCO = 1.0,
       tphlh$A$NCO = 1.0,
       tpllh$CI$S = 1.0,
       tplhl$CI$S = 1.0,
       tphlh$CI$S = 1.0,
       tphhl$CI$S = 1.0,
       tplhl$CI$NCO = 1.0,
       tphlh$CI$NCO = 1.0;

     // path delays
     (posedge CI *> (S +: !A)) = (tpllh$CI$S, tplhl$CI$S);
     (negedge CI *> (S +: A)) = (tphlh$CI$S, tphhl$CI$S);
     (CI *> NCO) = (tphlh$CI$NCO, tplhl$CI$NCO);
     (posedge A *> (S +: !CI)) = (tpllh$A$S, tplhl$A$S);
     (negedge A *> (S +: CI)) = (tphlh$A$S, tphhl$A$S);
     (A *> NCO) = (tphlh$A$NCO, tplhl$A$NCO);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_HA03D1 (CO, S, A, NCI);
input  A ;
input  NCI ;
output CO ;
output S ;

   not (I0_out, A);
   or  (I1_out, I0_out, NCI);
   not (CO, I1_out);
   xor (I3_out, A, NCI);
   not (S, I3_out);

   specify
     // delay parameters
     specparam
       tpllh$A$CO = 1.0,
       tphhl$A$CO = 1.0,
       tpllh$A$S = 1.0,
       tplhl$A$S = 1.0,
       tphlh$A$S = 1.0,
       tphhl$A$S = 1.0,
       tpllh$NCI$S = 1.0,
       tplhl$NCI$S = 1.0,
       tphlh$NCI$S = 1.0,
       tphhl$NCI$S = 1.0,
       tplhl$NCI$CO = 1.0,
       tphlh$NCI$CO = 1.0;

     // path delays
     (posedge NCI *> (S +: A)) = (tpllh$NCI$S, tplhl$NCI$S);
     (negedge NCI *> (S +: !A)) = (tphlh$NCI$S, tphhl$NCI$S);
     (NCI *> CO) = (tphlh$NCI$CO, tplhl$NCI$CO);
     (posedge A *> (S +: NCI)) = (tpllh$A$S, tplhl$A$S);
     (negedge A *> (S +: !NCI)) = (tphlh$A$S, tphhl$A$S);
     (A *> CO) = (tpllh$A$CO, tphhl$A$CO);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_HA03D2 (CO, S, A, NCI);
input  A ;
input  NCI ;
output CO ;
output S ;

   not (I0_out, A);
   or  (I1_out, I0_out, NCI);
   not (CO, I1_out);
   xor (I3_out, A, NCI);
   not (S, I3_out);

   specify
     // delay parameters
     specparam
       tpllh$A$CO = 1.0,
       tphhl$A$CO = 1.0,
       tpllh$A$S = 1.0,
       tplhl$A$S = 1.0,
       tphlh$A$S = 1.0,
       tphhl$A$S = 1.0,
       tpllh$NCI$S = 1.0,
       tplhl$NCI$S = 1.0,
       tphlh$NCI$S = 1.0,
       tphhl$NCI$S = 1.0,
       tplhl$NCI$CO = 1.0,
       tphlh$NCI$CO = 1.0;

     // path delays
     (posedge NCI *> (S +: A)) = (tpllh$NCI$S, tplhl$NCI$S);
     (negedge NCI *> (S +: !A)) = (tphlh$NCI$S, tphhl$NCI$S);
     (NCI *> CO) = (tphlh$NCI$CO, tplhl$NCI$CO);
     (posedge A *> (S +: NCI)) = (tpllh$A$S, tplhl$A$S);
     (negedge A *> (S +: !NCI)) = (tphlh$A$S, tphhl$A$S);
     (A *> CO) = (tpllh$A$CO, tphhl$A$CO);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_HA03D4 (CO, S, A, NCI);
input  A ;
input  NCI ;
output CO ;
output S ;

   not (I0_out, A);
   or  (I1_out, I0_out, NCI);
   not (CO, I1_out);
   xor (I3_out, A, NCI);
   not (S, I3_out);

   specify
     // delay parameters
     specparam
       tpllh$A$CO = 1.0,
       tphhl$A$CO = 1.0,
       tpllh$A$S = 1.0,
       tplhl$A$S = 1.0,
       tphlh$A$S = 1.0,
       tphhl$A$S = 1.0,
       tpllh$NCI$S = 1.0,
       tplhl$NCI$S = 1.0,
       tphlh$NCI$S = 1.0,
       tphhl$NCI$S = 1.0,
       tplhl$NCI$CO = 1.0,
       tphlh$NCI$CO = 1.0;

     // path delays
     (posedge NCI *> (S +: A)) = (tpllh$NCI$S, tplhl$NCI$S);
     (negedge NCI *> (S +: !A)) = (tphlh$NCI$S, tphhl$NCI$S);
     (NCI *> CO) = (tphlh$NCI$CO, tplhl$NCI$CO);
     (posedge A *> (S +: NCI)) = (tpllh$A$S, tplhl$A$S);
     (negedge A *> (S +: !NCI)) = (tphlh$A$S, tphhl$A$S);
     (A *> CO) = (tpllh$A$CO, tphhl$A$CO);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_IB01D12 (ZN, I);
input  I ;
output ZN ;

   not (ZN, I);

   specify
     // delay parameters
     specparam
       tplhl$I$ZN = 1.0,
       tphlh$I$ZN = 1.0;

     // path delays
     (I *> ZN) = (tphlh$I$ZN, tplhl$I$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_IB01D16 (ZN, I);
input  I ;
output ZN ;

   not (ZN, I);

   specify
     // delay parameters
     specparam
       tplhl$I$ZN = 1.0,
       tphlh$I$ZN = 1.0;

     // path delays
     (I *> ZN) = (tphlh$I$ZN, tplhl$I$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_IB01D8 (ZN, I);
input  I ;
output ZN ;

   not (ZN, I);

   specify
     // delay parameters
     specparam
       tplhl$I$ZN = 1.0,
       tphlh$I$ZN = 1.0;

     // path delays
     (I *> ZN) = (tphlh$I$ZN, tplhl$I$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_IN01D1 (ZN, I);
input  I ;
output ZN ;

   not (ZN, I);

   specify
     // delay parameters
     specparam
       tplhl$I$ZN = 1.0,
       tphlh$I$ZN = 1.0;

     // path delays
     (I *> ZN) = (tphlh$I$ZN, tplhl$I$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_IN01D12 (ZN, I);
input  I ;
output ZN ;

   not (ZN, I);

   specify
     // delay parameters
     specparam
       tplhl$I$ZN = 1.0,
       tphlh$I$ZN = 1.0;

     // path delays
     (I *> ZN) = (tphlh$I$ZN, tplhl$I$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_IN01D16 (ZN, I);
input  I ;
output ZN ;

   not (ZN, I);

   specify
     // delay parameters
     specparam
       tplhl$I$ZN = 1.0,
       tphlh$I$ZN = 1.0;

     // path delays
     (I *> ZN) = (tphlh$I$ZN, tplhl$I$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_IN01D2 (ZN, I);
input  I ;
output ZN ;

   not (ZN, I);

   specify
     // delay parameters
     specparam
       tplhl$I$ZN = 1.0,
       tphlh$I$ZN = 1.0;

     // path delays
     (I *> ZN) = (tphlh$I$ZN, tplhl$I$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_IN01D3 (ZN, I);
input  I ;
output ZN ;

   not (ZN, I);

   specify
     // delay parameters
     specparam
       tplhl$I$ZN = 1.0,
       tphlh$I$ZN = 1.0;

     // path delays
     (I *> ZN) = (tphlh$I$ZN, tplhl$I$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_IN01D4 (ZN, I);
input  I ;
output ZN ;

   not (ZN, I);

   specify
     // delay parameters
     specparam
       tplhl$I$ZN = 1.0,
       tphlh$I$ZN = 1.0;

     // path delays
     (I *> ZN) = (tphlh$I$ZN, tplhl$I$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_IN01D6 (ZN, I);
input  I ;
output ZN ;

   not (ZN, I);

   specify
     // delay parameters
     specparam
       tplhl$I$ZN = 1.0,
       tphlh$I$ZN = 1.0;

     // path delays
     (I *> ZN) = (tphlh$I$ZN, tplhl$I$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_IN01D8 (ZN, I);
input  I ;
output ZN ;

   not (ZN, I);

   specify
     // delay parameters
     specparam
       tplhl$I$ZN = 1.0,
       tphlh$I$ZN = 1.0;

     // path delays
     (I *> ZN) = (tphlh$I$ZN, tplhl$I$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_IT01D1 (ZN, I, OE);
input  I ;
input  OE ;
output ZN ;

   not (I0_out, I);
   bufif1 (ZN, I0_out, OE);

   specify
     // delay parameters
     specparam
       tplhl$I$ZN = 1.0,
       tphlh$I$ZN = 1.0,
       tpzh$OE$ZN = 1.0,
       tpzl$OE$ZN = 1.0,
       tplz$OE$ZN = 1.0,
       tphz$OE$ZN = 1.0;

     // path delays
     (OE *> ZN) = (0, 0, tplz$OE$ZN, tpzh$OE$ZN, tphz$OE$ZN, tpzl$OE$ZN);
     (I *> ZN) = (tphlh$I$ZN, tplhl$I$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_IT01D2 (ZN, I, OE);
input  I ;
input  OE ;
output ZN ;

   not (I0_out, I);
   bufif1 (ZN, I0_out, OE);

   specify
     // delay parameters
     specparam
       tplhl$I$ZN = 1.0,
       tphlh$I$ZN = 1.0,
       tpzh$OE$ZN = 1.0,
       tpzl$OE$ZN = 1.0,
       tplz$OE$ZN = 1.0,
       tphz$OE$ZN = 1.0;

     // path delays
     (OE *> ZN) = (0, 0, tplz$OE$ZN, tpzh$OE$ZN, tphz$OE$ZN, tpzl$OE$ZN);
     (I *> ZN) = (tphlh$I$ZN, tplhl$I$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_IT01D4 (ZN, I, OE);
input  I ;
input  OE ;
output ZN ;

   not (I0_out, I);
   bufif1 (ZN, I0_out, OE);

   specify
     // delay parameters
     specparam
       tplhl$I$ZN = 1.0,
       tphlh$I$ZN = 1.0,
       tpzh$OE$ZN = 1.0,
       tpzl$OE$ZN = 1.0,
       tplz$OE$ZN = 1.0,
       tphz$OE$ZN = 1.0;

     // path delays
     (OE *> ZN) = (0, 0, tplz$OE$ZN, tpzh$OE$ZN, tphz$OE$ZN, tpzl$OE$ZN);
     (I *> ZN) = (tphlh$I$ZN, tplhl$I$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_IT01D6 (ZN, I, OE);
input  I ;
input  OE ;
output ZN ;

   not (I0_out, I);
   bufif1 (ZN, I0_out, OE);

   specify
     // delay parameters
     specparam
       tplhl$I$ZN = 1.0,
       tphlh$I$ZN = 1.0,
       tpzh$OE$ZN = 1.0,
       tpzl$OE$ZN = 1.0,
       tplz$OE$ZN = 1.0,
       tphz$OE$ZN = 1.0;

     // path delays
     (OE *> ZN) = (0, 0, tplz$OE$ZN, tpzh$OE$ZN, tphz$OE$ZN, tpzl$OE$ZN);
     (I *> ZN) = (tphlh$I$ZN, tplhl$I$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_IT02D1 (ZN, I, OE);
input  I ;
input  OE ;
output ZN ;

   not (I0_out, I);
   bufif0 (ZN, I0_out, OE);

   specify
     // delay parameters
     specparam
       tplhl$I$ZN = 1.0,
       tphlh$I$ZN = 1.0,
       tplz$OE$ZN = 1.0,
       tphz$OE$ZN = 1.0,
       tpzh$OE$ZN = 1.0,
       tpzl$OE$ZN = 1.0;

     // path delays
     (OE *> ZN) = (0, 0, tplz$OE$ZN, tpzh$OE$ZN, tphz$OE$ZN, tpzl$OE$ZN);
     (I *> ZN) = (tphlh$I$ZN, tplhl$I$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_IT02D2 (ZN, I, OE);
input  I ;
input  OE ;
output ZN ;

   not (I0_out, I);
   bufif0 (ZN, I0_out, OE);

   specify
     // delay parameters
     specparam
       tplhl$I$ZN = 1.0,
       tphlh$I$ZN = 1.0,
       tplz$OE$ZN = 1.0,
       tphz$OE$ZN = 1.0,
       tpzh$OE$ZN = 1.0,
       tpzl$OE$ZN = 1.0;

     // path delays
     (OE *> ZN) = (0, 0, tplz$OE$ZN, tpzh$OE$ZN, tphz$OE$ZN, tpzl$OE$ZN);
     (I *> ZN) = (tphlh$I$ZN, tplhl$I$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_IT02D4 (ZN, I, OE);
input  I ;
input  OE ;
output ZN ;

   not (I0_out, I);
   bufif0 (ZN, I0_out, OE);

   specify
     // delay parameters
     specparam
       tplhl$I$ZN = 1.0,
       tphlh$I$ZN = 1.0,
       tplz$OE$ZN = 1.0,
       tphz$OE$ZN = 1.0,
       tpzh$OE$ZN = 1.0,
       tpzl$OE$ZN = 1.0;

     // path delays
     (OE *> ZN) = (0, 0, tplz$OE$ZN, tpzh$OE$ZN, tphz$OE$ZN, tpzl$OE$ZN);
     (I *> ZN) = (tphlh$I$ZN, tplhl$I$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_IT02D6 (ZN, I, OE);
input  I ;
input  OE ;
output ZN ;

   not (I0_out, I);
   bufif0 (ZN, I0_out, OE);

   specify
     // delay parameters
     specparam
       tplhl$I$ZN = 1.0,
       tphlh$I$ZN = 1.0,
       tplz$OE$ZN = 1.0,
       tphz$OE$ZN = 1.0,
       tpzh$OE$ZN = 1.0,
       tpzl$OE$ZN = 1.0;

     // path delays
     (OE *> ZN) = (0, 0, tplz$OE$ZN, tpzh$OE$ZN, tphz$OE$ZN, tpzl$OE$ZN);
     (I *> ZN) = (tphlh$I$ZN, tplhl$I$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_MA01D1 (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   and (I0_out, A, B);
   and (I1_out, B, C);
   and (I3_out, C, A);
   or  (Z, I0_out, I1_out, I3_out);

   specify
     // delay parameters
     specparam
       tpllh$A$Z = 1.0,
       tphhl$A$Z = 1.0,
       tpllh$B$Z = 1.0,
       tphhl$B$Z = 1.0,
       tpllh$C$Z = 1.0,
       tphhl$C$Z = 1.0,
       tpllh$A$Z$B_EQ_0_AN_C_EQ_1 = 1.0,
       tphhl$A$Z$B_EQ_0_AN_C_EQ_1 = 1.0,
       tpllh$A$Z$B_EQ_1_AN_C_EQ_0 = 1.0,
       tphhl$A$Z$B_EQ_1_AN_C_EQ_0 = 1.0,
       tpllh$B$Z$A_EQ_1_AN_C_EQ_0 = 1.0,
       tphhl$B$Z$A_EQ_1_AN_C_EQ_0 = 1.0,
       tpllh$B$Z$A_EQ_0_AN_C_EQ_1 = 1.0,
       tphhl$B$Z$A_EQ_0_AN_C_EQ_1 = 1.0,
       tpllh$C$Z$A_EQ_0_AN_B_EQ_1 = 1.0,
       tphhl$C$Z$A_EQ_0_AN_B_EQ_1 = 1.0,
       tpllh$C$Z$A_EQ_1_AN_B_EQ_0 = 1.0,
       tphhl$C$Z$A_EQ_1_AN_B_EQ_0 = 1.0;

     // path delays
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (tpllh$C$Z$A_EQ_1_AN_B_EQ_0, tphhl$C$Z$A_EQ_1_AN_B_EQ_0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (tpllh$C$Z$A_EQ_0_AN_B_EQ_1, tphhl$C$Z$A_EQ_0_AN_B_EQ_1);
     ifnone
       (C *> Z) = (tpllh$C$Z,tphhl$C$Z);

     if (A == 1'b1 && C == 1'b0)
       (B *> Z) = (tpllh$B$Z$A_EQ_1_AN_C_EQ_0, tphhl$B$Z$A_EQ_1_AN_C_EQ_0);
     if (A == 1'b0 && C == 1'b1)
       (B *> Z) = (tpllh$B$Z$A_EQ_0_AN_C_EQ_1, tphhl$B$Z$A_EQ_0_AN_C_EQ_1);
     ifnone
       (B *> Z) = (tpllh$B$Z,tphhl$B$Z);

     if (B == 1'b1 && C == 1'b0)
       (A *> Z) = (tpllh$A$Z$B_EQ_1_AN_C_EQ_0, tphhl$A$Z$B_EQ_1_AN_C_EQ_0);
     if (B == 1'b0 && C == 1'b1)
       (A *> Z) = (tpllh$A$Z$B_EQ_0_AN_C_EQ_1, tphhl$A$Z$B_EQ_0_AN_C_EQ_1);
     ifnone
       (A *> Z) = (tpllh$A$Z,tphhl$A$Z);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_MA01D2 (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   and (I0_out, A, B);
   and (I1_out, B, C);
   and (I3_out, C, A);
   or  (Z, I0_out, I1_out, I3_out);

   specify
     // delay parameters
     specparam
       tpllh$A$Z = 1.0,
       tphhl$A$Z = 1.0,
       tpllh$B$Z = 1.0,
       tphhl$B$Z = 1.0,
       tpllh$C$Z = 1.0,
       tphhl$C$Z = 1.0,
       tpllh$A$Z$B_EQ_0_AN_C_EQ_1 = 1.0,
       tphhl$A$Z$B_EQ_0_AN_C_EQ_1 = 1.0,
       tpllh$A$Z$B_EQ_1_AN_C_EQ_0 = 1.0,
       tphhl$A$Z$B_EQ_1_AN_C_EQ_0 = 1.0,
       tpllh$B$Z$A_EQ_1_AN_C_EQ_0 = 1.0,
       tphhl$B$Z$A_EQ_1_AN_C_EQ_0 = 1.0,
       tpllh$B$Z$A_EQ_0_AN_C_EQ_1 = 1.0,
       tphhl$B$Z$A_EQ_0_AN_C_EQ_1 = 1.0,
       tpllh$C$Z$A_EQ_0_AN_B_EQ_1 = 1.0,
       tphhl$C$Z$A_EQ_0_AN_B_EQ_1 = 1.0,
       tpllh$C$Z$A_EQ_1_AN_B_EQ_0 = 1.0,
       tphhl$C$Z$A_EQ_1_AN_B_EQ_0 = 1.0;

     // path delays
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (tpllh$C$Z$A_EQ_1_AN_B_EQ_0, tphhl$C$Z$A_EQ_1_AN_B_EQ_0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (tpllh$C$Z$A_EQ_0_AN_B_EQ_1, tphhl$C$Z$A_EQ_0_AN_B_EQ_1);
     ifnone
       (C *> Z) = (tpllh$C$Z,tphhl$C$Z);

     if (A == 1'b1 && C == 1'b0)
       (B *> Z) = (tpllh$B$Z$A_EQ_1_AN_C_EQ_0, tphhl$B$Z$A_EQ_1_AN_C_EQ_0);
     if (A == 1'b0 && C == 1'b1)
       (B *> Z) = (tpllh$B$Z$A_EQ_0_AN_C_EQ_1, tphhl$B$Z$A_EQ_0_AN_C_EQ_1);
     ifnone
       (B *> Z) = (tpllh$B$Z,tphhl$B$Z);

     if (B == 1'b1 && C == 1'b0)
       (A *> Z) = (tpllh$A$Z$B_EQ_1_AN_C_EQ_0, tphhl$A$Z$B_EQ_1_AN_C_EQ_0);
     if (B == 1'b0 && C == 1'b1)
       (A *> Z) = (tpllh$A$Z$B_EQ_0_AN_C_EQ_1, tphhl$A$Z$B_EQ_0_AN_C_EQ_1);
     ifnone
       (A *> Z) = (tpllh$A$Z,tphhl$A$Z);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_MA01D4 (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   and (I0_out, A, B);
   and (I1_out, B, C);
   and (I3_out, C, A);
   or  (Z, I0_out, I1_out, I3_out);

   specify
     // delay parameters
     specparam
       tpllh$A$Z = 1.0,
       tphhl$A$Z = 1.0,
       tpllh$B$Z = 1.0,
       tphhl$B$Z = 1.0,
       tpllh$C$Z = 1.0,
       tphhl$C$Z = 1.0,
       tpllh$A$Z$B_EQ_0_AN_C_EQ_1 = 1.0,
       tphhl$A$Z$B_EQ_0_AN_C_EQ_1 = 1.0,
       tpllh$A$Z$B_EQ_1_AN_C_EQ_0 = 1.0,
       tphhl$A$Z$B_EQ_1_AN_C_EQ_0 = 1.0,
       tpllh$B$Z$A_EQ_1_AN_C_EQ_0 = 1.0,
       tphhl$B$Z$A_EQ_1_AN_C_EQ_0 = 1.0,
       tpllh$B$Z$A_EQ_0_AN_C_EQ_1 = 1.0,
       tphhl$B$Z$A_EQ_0_AN_C_EQ_1 = 1.0,
       tpllh$C$Z$A_EQ_0_AN_B_EQ_1 = 1.0,
       tphhl$C$Z$A_EQ_0_AN_B_EQ_1 = 1.0,
       tpllh$C$Z$A_EQ_1_AN_B_EQ_0 = 1.0,
       tphhl$C$Z$A_EQ_1_AN_B_EQ_0 = 1.0;

     // path delays
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (tpllh$C$Z$A_EQ_1_AN_B_EQ_0, tphhl$C$Z$A_EQ_1_AN_B_EQ_0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (tpllh$C$Z$A_EQ_0_AN_B_EQ_1, tphhl$C$Z$A_EQ_0_AN_B_EQ_1);
     ifnone
       (C *> Z) = (tpllh$C$Z,tphhl$C$Z);

     if (A == 1'b1 && C == 1'b0)
       (B *> Z) = (tpllh$B$Z$A_EQ_1_AN_C_EQ_0, tphhl$B$Z$A_EQ_1_AN_C_EQ_0);
     if (A == 1'b0 && C == 1'b1)
       (B *> Z) = (tpllh$B$Z$A_EQ_0_AN_C_EQ_1, tphhl$B$Z$A_EQ_0_AN_C_EQ_1);
     ifnone
       (B *> Z) = (tpllh$B$Z,tphhl$B$Z);

     if (B == 1'b1 && C == 1'b0)
       (A *> Z) = (tpllh$A$Z$B_EQ_1_AN_C_EQ_0, tphhl$A$Z$B_EQ_1_AN_C_EQ_0);
     if (B == 1'b0 && C == 1'b1)
       (A *> Z) = (tpllh$A$Z$B_EQ_0_AN_C_EQ_1, tphhl$A$Z$B_EQ_0_AN_C_EQ_1);
     ifnone
       (A *> Z) = (tpllh$A$Z,tphhl$A$Z);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_MX02D1 (Z, I0, I1, OE);
input  I0 ;
input  I1 ;
input  OE ;
output Z ;

   udp_mux2 (Z, I0, I1, OE);

   specify
     // delay parameters
     specparam
       tpllh$I0$Z = 1.0,
       tphhl$I0$Z = 1.0,
       tpllh$I1$Z = 1.0,
       tphhl$I1$Z = 1.0,
       tpllh$OE$Z = 1.0,
       tplhl$OE$Z = 1.0,
       tphlh$OE$Z = 1.0,
       tphhl$OE$Z = 1.0,
       tpllh$I0$Z$I1_EQ_1_AN_OE_EQ_0 = 1.0,
       tphhl$I0$Z$I1_EQ_1_AN_OE_EQ_0 = 1.0,
       tpllh$I0$Z$I1_EQ_0_AN_OE_EQ_0 = 1.0,
       tphhl$I0$Z$I1_EQ_0_AN_OE_EQ_0 = 1.0,
       tpllh$I1$Z$I0_EQ_1_AN_OE_EQ_1 = 1.0,
       tphhl$I1$Z$I0_EQ_1_AN_OE_EQ_1 = 1.0,
       tpllh$I1$Z$I0_EQ_0_AN_OE_EQ_1 = 1.0,
       tphhl$I1$Z$I0_EQ_0_AN_OE_EQ_1 = 1.0;

     // path delays
     (posedge OE *> (Z +: I1)) = (tpllh$OE$Z, tplhl$OE$Z);
     (negedge OE *> (Z +: I0)) = (tphlh$OE$Z, tphhl$OE$Z);
     if (I0 == 1'b1 && OE == 1'b1)
       (I1 *> Z) = (tpllh$I1$Z$I0_EQ_1_AN_OE_EQ_1, tphhl$I1$Z$I0_EQ_1_AN_OE_EQ_1);
     if (I0 == 1'b0 && OE == 1'b1)
       (I1 *> Z) = (tpllh$I1$Z$I0_EQ_0_AN_OE_EQ_1, tphhl$I1$Z$I0_EQ_0_AN_OE_EQ_1);
     ifnone
       (I1 *> Z) = (tpllh$I1$Z,tphhl$I1$Z);

     if (I1 == 1'b1 && OE == 1'b0)
       (I0 *> Z) = (tpllh$I0$Z$I1_EQ_1_AN_OE_EQ_0, tphhl$I0$Z$I1_EQ_1_AN_OE_EQ_0);
     if (I1 == 1'b0 && OE == 1'b0)
       (I0 *> Z) = (tpllh$I0$Z$I1_EQ_0_AN_OE_EQ_0, tphhl$I0$Z$I1_EQ_0_AN_OE_EQ_0);
     ifnone
       (I0 *> Z) = (tpllh$I0$Z,tphhl$I0$Z);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_MX02D2 (Z, I0, I1, OE);
input  I0 ;
input  I1 ;
input  OE ;
output Z ;

   udp_mux2 (Z, I0, I1, OE);

   specify
     // delay parameters
     specparam
       tpllh$I0$Z = 1.0,
       tphhl$I0$Z = 1.0,
       tpllh$I1$Z = 1.0,
       tphhl$I1$Z = 1.0,
       tpllh$OE$Z = 1.0,
       tplhl$OE$Z = 1.0,
       tphlh$OE$Z = 1.0,
       tphhl$OE$Z = 1.0,
       tpllh$I0$Z$I1_EQ_1_AN_OE_EQ_0 = 1.0,
       tphhl$I0$Z$I1_EQ_1_AN_OE_EQ_0 = 1.0,
       tpllh$I0$Z$I1_EQ_0_AN_OE_EQ_0 = 1.0,
       tphhl$I0$Z$I1_EQ_0_AN_OE_EQ_0 = 1.0,
       tpllh$I1$Z$I0_EQ_0_AN_OE_EQ_1 = 1.0,
       tphhl$I1$Z$I0_EQ_0_AN_OE_EQ_1 = 1.0,
       tpllh$I1$Z$I0_EQ_1_AN_OE_EQ_1 = 1.0,
       tphhl$I1$Z$I0_EQ_1_AN_OE_EQ_1 = 1.0;

     // path delays
     (posedge OE *> (Z +: I1)) = (tpllh$OE$Z, tplhl$OE$Z);
     (negedge OE *> (Z +: I0)) = (tphlh$OE$Z, tphhl$OE$Z);
     if (I0 == 1'b1 && OE == 1'b1)
       (I1 *> Z) = (tpllh$I1$Z$I0_EQ_1_AN_OE_EQ_1, tphhl$I1$Z$I0_EQ_1_AN_OE_EQ_1);
     if (I0 == 1'b0 && OE == 1'b1)
       (I1 *> Z) = (tpllh$I1$Z$I0_EQ_0_AN_OE_EQ_1, tphhl$I1$Z$I0_EQ_0_AN_OE_EQ_1);
     ifnone
       (I1 *> Z) = (tpllh$I1$Z,tphhl$I1$Z);

     if (I1 == 1'b1 && OE == 1'b0)
       (I0 *> Z) = (tpllh$I0$Z$I1_EQ_1_AN_OE_EQ_0, tphhl$I0$Z$I1_EQ_1_AN_OE_EQ_0);
     if (I1 == 1'b0 && OE == 1'b0)
       (I0 *> Z) = (tpllh$I0$Z$I1_EQ_0_AN_OE_EQ_0, tphhl$I0$Z$I1_EQ_0_AN_OE_EQ_0);
     ifnone
       (I0 *> Z) = (tpllh$I0$Z,tphhl$I0$Z);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_MX02D4 (Z, I0, I1, OE);
input  I0 ;
input  I1 ;
input  OE ;
output Z ;

   udp_mux2 (Z, I0, I1, OE);

   specify
     // delay parameters
     specparam
       tpllh$I0$Z = 1.0,
       tphhl$I0$Z = 1.0,
       tpllh$I1$Z = 1.0,
       tphhl$I1$Z = 1.0,
       tpllh$OE$Z = 1.0,
       tplhl$OE$Z = 1.0,
       tphlh$OE$Z = 1.0,
       tphhl$OE$Z = 1.0,
       tpllh$I0$Z$I1_EQ_1_AN_OE_EQ_0 = 1.0,
       tphhl$I0$Z$I1_EQ_1_AN_OE_EQ_0 = 1.0,
       tpllh$I0$Z$I1_EQ_0_AN_OE_EQ_0 = 1.0,
       tphhl$I0$Z$I1_EQ_0_AN_OE_EQ_0 = 1.0,
       tpllh$I1$Z$I0_EQ_0_AN_OE_EQ_1 = 1.0,
       tphhl$I1$Z$I0_EQ_0_AN_OE_EQ_1 = 1.0,
       tpllh$I1$Z$I0_EQ_1_AN_OE_EQ_1 = 1.0,
       tphhl$I1$Z$I0_EQ_1_AN_OE_EQ_1 = 1.0;

     // path delays
     (posedge OE *> (Z +: I1)) = (tpllh$OE$Z, tplhl$OE$Z);
     (negedge OE *> (Z +: I0)) = (tphlh$OE$Z, tphhl$OE$Z);
     if (I0 == 1'b1 && OE == 1'b1)
       (I1 *> Z) = (tpllh$I1$Z$I0_EQ_1_AN_OE_EQ_1, tphhl$I1$Z$I0_EQ_1_AN_OE_EQ_1);
     if (I0 == 1'b0 && OE == 1'b1)
       (I1 *> Z) = (tpllh$I1$Z$I0_EQ_0_AN_OE_EQ_1, tphhl$I1$Z$I0_EQ_0_AN_OE_EQ_1);
     ifnone
       (I1 *> Z) = (tpllh$I1$Z,tphhl$I1$Z);

     if (I1 == 1'b1 && OE == 1'b0)
       (I0 *> Z) = (tpllh$I0$Z$I1_EQ_1_AN_OE_EQ_0, tphhl$I0$Z$I1_EQ_1_AN_OE_EQ_0);
     if (I1 == 1'b0 && OE == 1'b0)
       (I0 *> Z) = (tpllh$I0$Z$I1_EQ_0_AN_OE_EQ_0, tphhl$I0$Z$I1_EQ_0_AN_OE_EQ_0);
     ifnone
       (I0 *> Z) = (tpllh$I0$Z,tphhl$I0$Z);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_MX03D1 (Z, I0, I1, I2, OE0, OE1);
input  I0 ;
input  I1 ;
input  I2 ;
input  OE0 ;
input  OE1 ;
output Z ;

   udp_mux2 (I0_out, I0, I1, OE0);
   udp_mux2 (Z, I0_out, I2, OE1);

   specify
     // delay parameters
     specparam
       tpllh$I0$Z = 1.0,
       tphhl$I0$Z = 1.0,
       tpllh$I1$Z = 1.0,
       tphhl$I1$Z = 1.0,
       tpllh$I2$Z = 1.0,
       tphhl$I2$Z = 1.0,
       tpllh$OE0$Z = 1.0,
       tplhl$OE0$Z = 1.0,
       tphlh$OE0$Z = 1.0,
       tphhl$OE0$Z = 1.0,
       tpllh$OE1$Z = 1.0,
       tplhl$OE1$Z = 1.0,
       tphlh$OE1$Z = 1.0,
       tphhl$OE1$Z = 1.0,
       tpllh$I0$Z$I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphhl$I0$Z$I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tpllh$I0$Z$I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphhl$I0$Z$I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tpllh$I1$Z$I0_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tphhl$I1$Z$I0_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tpllh$I1$Z$I0_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tphhl$I1$Z$I0_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tpllh$I2$Z$I0_EQ_1_AN_I1_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1 = 1.0,
       tphhl$I2$Z$I0_EQ_1_AN_I1_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1 = 1.0,
       tpllh$I2$Z$I0_EQ_0_AN_I1_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1 = 1.0,
       tphhl$I2$Z$I0_EQ_0_AN_I1_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1 = 1.0,
       tpllh$OE0$Z$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphhl$OE0$Z$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE1_EQ_0 = 1.0,
       tpllh$OE0$Z$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE1_EQ_0 = 1.0,
       tphhl$OE0$Z$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE1_EQ_0 = 1.0,
       tplhl$OE0$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphlh$OE0$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE1_EQ_0 = 1.0,
       tplhl$OE0$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE1_EQ_0 = 1.0,
       tphlh$OE0$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE1_EQ_0 = 1.0,
       tpllh$OE1$Z$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_0 = 1.0,
       tphhl$OE1$Z$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_0 = 1.0,
       tpllh$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_1 = 1.0,
       tphhl$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_1 = 1.0,
       tplhl$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0 = 1.0,
       tphlh$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0 = 1.0,
       tplhl$OE1$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE0_EQ_1 = 1.0,
       tphlh$OE1$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE0_EQ_1 = 1.0;

     // path delays
      (posedge OE1 => (Z +: Z)) = (1.0, 1.0);
      (negedge OE1 => (Z -: Z)) = (1.0, 1.0);

     if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && OE0 == 1'b1)
       (OE1 *> Z) = (tphlh$OE1$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE0_EQ_1, tplhl$OE1$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE0_EQ_1);
     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && OE0 == 1'b1)
       (OE1 *> Z) = (tpllh$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_1, tphhl$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_1);
     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && OE0 == 1'b0)
       (OE1 *> Z) = (tphlh$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0, tplhl$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0);
     if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && OE0 == 1'b0)
       (OE1 *> Z) = (tpllh$OE1$Z$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_0, tphhl$OE1$Z$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_0);
  //   ifnone
   //    (OE1 *> Z) = (tpllh$OE1$Z,tplhl$OE1$Z);

      (posedge OE0 => (Z +: Z)) = (1.0, 1.0);
      (negedge OE0 => (Z -: Z)) = (1.0, 1.0);

     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && OE1 == 1'b0)
       (OE0 *> Z) = (tphlh$OE0$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE1_EQ_0, tplhl$OE0$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE1_EQ_0);
     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && OE1 == 1'b0)
       (OE0 *> Z) = (tphlh$OE0$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE1_EQ_0, tplhl$OE0$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE1_EQ_0);
     if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && OE1 == 1'b0)
       (OE0 *> Z) = (tpllh$OE0$Z$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE1_EQ_0, tphhl$OE0$Z$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE1_EQ_0);
     if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && OE1 == 1'b0)
       (OE0 *> Z) = (tpllh$OE0$Z$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE1_EQ_0, tphhl$OE0$Z$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE1_EQ_0);
    // ifnone
     //  (OE0 *> Z) = (tpllh$OE0$Z,tplhl$OE0$Z);
      (posedge I2 => (Z +: Z)) = (1.0, 1.0);
     if (I0 == 1'b1 && I1 == 1'b1 && OE0 == 1'b1 && OE1 == 1'b1)
       (I2 *> Z) = (tpllh$I2$Z$I0_EQ_1_AN_I1_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1, tphhl$I2$Z$I0_EQ_1_AN_I1_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1);
     if (I0 == 1'b0 && I1 == 1'b0 && OE0 == 1'b0 && OE1 == 1'b1)
       (I2 *> Z) = (tpllh$I2$Z$I0_EQ_0_AN_I1_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1, tphhl$I2$Z$I0_EQ_0_AN_I1_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1);
    // ifnone
 //      (I2 *> Z) = (tpllh$I2$Z,tphhl$I2$Z);
      (posedge I1 => (Z +: Z)) = (1.0, 1.0);
     if (I0 == 1'b1 && I2 == 1'b1 && OE0 == 1'b1 && OE1 == 1'b0)
       (I1 *> Z) = (tpllh$I1$Z$I0_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0, tphhl$I1$Z$I0_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0);
     if (I0 == 1'b0 && I2 == 1'b0 && OE0 == 1'b1 && OE1 == 1'b0)
       (I1 *> Z) = (tpllh$I1$Z$I0_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0, tphhl$I1$Z$I0_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0);
   //  ifnone
   //    (I1 *> Z) = (tpllh$I1$Z,tphhl$I1$Z);
      (posedge I0 => (Z +: Z)) = (1.0, 1.0);
     if (I1 == 1'b1 && I2 == 1'b1 && OE0 == 1'b0 && OE1 == 1'b0)
       (I0 *> Z) = (tpllh$I0$Z$I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0, tphhl$I0$Z$I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0);
     if (I1 == 1'b0 && I2 == 1'b0 && OE0 == 1'b0 && OE1 == 1'b0)
       (I0 *> Z) = (tpllh$I0$Z$I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0, tphhl$I0$Z$I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0);
  //   ifnone
  //     (I0 *> Z) = (tpllh$I0$Z,tphhl$I0$Z);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_MX03D2 (Z, I0, I1, I2, OE0, OE1);
input  I0 ;
input  I1 ;
input  I2 ;
input  OE0 ;
input  OE1 ;
output Z ;

   udp_mux2 (I0_out, I0, I1, OE0);
   udp_mux2 (Z, I0_out, I2, OE1);

   specify
     // delay parameters
     specparam
       tpllh$I0$Z = 1.0,
       tphhl$I0$Z = 1.0,
       tpllh$I1$Z = 1.0,
       tphhl$I1$Z = 1.0,
       tpllh$I2$Z = 1.0,
       tphhl$I2$Z = 1.0,
       tpllh$OE0$Z = 1.0,
       tplhl$OE0$Z = 1.0,
       tphlh$OE0$Z = 1.0,
       tphhl$OE0$Z = 1.0,
       tpllh$OE1$Z = 1.0,
       tplhl$OE1$Z = 1.0,
       tphlh$OE1$Z = 1.0,
       tphhl$OE1$Z = 1.0,
       tpllh$I0$Z$I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphhl$I0$Z$I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tpllh$I0$Z$I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphhl$I0$Z$I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tpllh$I1$Z$I0_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tphhl$I1$Z$I0_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tpllh$I1$Z$I0_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tphhl$I1$Z$I0_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tpllh$I2$Z$I0_EQ_0_AN_I1_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1 = 1.0,
       tphhl$I2$Z$I0_EQ_0_AN_I1_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1 = 1.0,
       tpllh$I2$Z$I0_EQ_1_AN_I1_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1 = 1.0,
       tphhl$I2$Z$I0_EQ_1_AN_I1_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1 = 1.0,
       tpllh$OE0$Z$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphhl$OE0$Z$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE1_EQ_0 = 1.0,
       tpllh$OE0$Z$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE1_EQ_0 = 1.0,
       tphhl$OE0$Z$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE1_EQ_0 = 1.0,
       tplhl$OE0$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphlh$OE0$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE1_EQ_0 = 1.0,
       tplhl$OE0$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE1_EQ_0 = 1.0,
       tphlh$OE0$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE1_EQ_0 = 1.0,
       tpllh$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_1 = 1.0,
       tphhl$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_1 = 1.0,
       tpllh$OE1$Z$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_0 = 1.0,
       tphhl$OE1$Z$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_0 = 1.0,
       tplhl$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0 = 1.0,
       tphlh$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0 = 1.0,
       tplhl$OE1$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE0_EQ_1 = 1.0,
       tphlh$OE1$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE0_EQ_1 = 1.0;

     // path delays

      (posedge OE1 => (Z +: Z)) = (1.0, 1.0);
      (negedge OE1 => (Z -: Z)) = (1.0, 1.0);
     if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && OE0 == 1'b1)
       (OE1 *> Z) = (tphlh$OE1$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE0_EQ_1, tplhl$OE1$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE0_EQ_1);
     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && OE0 == 1'b1)
       (OE1 *> Z) = (tpllh$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_1, tphhl$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_1);
     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && OE0 == 1'b0)
       (OE1 *> Z) = (tphlh$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0, tplhl$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0);
     if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && OE0 == 1'b0)
       (OE1 *> Z) = (tpllh$OE1$Z$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_0, tphhl$OE1$Z$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_0);
   //  ifnone
  //     (OE1 *> Z) = (tpllh$OE1$Z,tplhl$OE1$Z);

      (posedge OE0 => (Z +: Z)) = (1.0, 1.0);
      (negedge OE0 => (Z -: Z)) = (1.0, 1.0);
     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && OE1 == 1'b0)
       (OE0 *> Z) = (tphlh$OE0$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE1_EQ_0, tplhl$OE0$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE1_EQ_0);
     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && OE1 == 1'b0)
       (OE0 *> Z) = (tphlh$OE0$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE1_EQ_0, tplhl$OE0$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE1_EQ_0);
     if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && OE1 == 1'b0)
       (OE0 *> Z) = (tpllh$OE0$Z$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE1_EQ_0, tphhl$OE0$Z$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE1_EQ_0);
     if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && OE1 == 1'b0)
       (OE0 *> Z) = (tpllh$OE0$Z$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE1_EQ_0, tphhl$OE0$Z$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE1_EQ_0);
//     ifnone
   //    (OE0 *> Z) = (tpllh$OE0$Z,tplhl$OE0$Z);

      (posedge I2 => (Z +: Z)) = (1.0, 1.0);
     if (I0 == 1'b1 && I1 == 1'b1 && OE0 == 1'b1 && OE1 == 1'b1)
       (I2 *> Z) = (tpllh$I2$Z$I0_EQ_1_AN_I1_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1, tphhl$I2$Z$I0_EQ_1_AN_I1_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1);
     if (I0 == 1'b0 && I1 == 1'b0 && OE0 == 1'b0 && OE1 == 1'b1)
       (I2 *> Z) = (tpllh$I2$Z$I0_EQ_0_AN_I1_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1, tphhl$I2$Z$I0_EQ_0_AN_I1_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1);
    // ifnone
    //   (I2 *> Z) = (tpllh$I2$Z,tphhl$I2$Z);

      (posedge I1 => (Z +: Z)) = (1.0, 1.0);
     if (I0 == 1'b1 && I2 == 1'b1 && OE0 == 1'b1 && OE1 == 1'b0)
       (I1 *> Z) = (tpllh$I1$Z$I0_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0, tphhl$I1$Z$I0_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0);
     if (I0 == 1'b0 && I2 == 1'b0 && OE0 == 1'b1 && OE1 == 1'b0)
       (I1 *> Z) = (tpllh$I1$Z$I0_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0, tphhl$I1$Z$I0_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0);
  //   ifnone
   //    (I1 *> Z) = (tpllh$I1$Z,tphhl$I1$Z);
      (posedge I0 => (Z +: Z)) = (1.0, 1.0);
     if (I1 == 1'b1 && I2 == 1'b1 && OE0 == 1'b0 && OE1 == 1'b0)
       (I0 *> Z) = (tpllh$I0$Z$I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0, tphhl$I0$Z$I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0);
     if (I1 == 1'b0 && I2 == 1'b0 && OE0 == 1'b0 && OE1 == 1'b0)
       (I0 *> Z) = (tpllh$I0$Z$I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0, tphhl$I0$Z$I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0);
  //   ifnone
  //     (I0 *> Z) = (tpllh$I0$Z,tphhl$I0$Z);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_MX03D4 (Z, I0, I1, I2, OE0, OE1);
input  I0 ;
input  I1 ;
input  I2 ;
input  OE0 ;
input  OE1 ;
output Z ;

   udp_mux2 (I0_out, I0, I1, OE0);
   udp_mux2 (Z, I0_out, I2, OE1);

   specify
     // delay parameters
     specparam
       tpllh$I0$Z = 1.0,
       tphhl$I0$Z = 1.0,
       tpllh$I1$Z = 1.0,
       tphhl$I1$Z = 1.0,
       tpllh$I2$Z = 1.0,
       tphhl$I2$Z = 1.0,
       tpllh$OE0$Z = 1.0,
       tplhl$OE0$Z = 1.0,
       tphlh$OE0$Z = 1.0,
       tphhl$OE0$Z = 1.0,
       tpllh$OE1$Z = 1.0,
       tplhl$OE1$Z = 1.0,
       tphlh$OE1$Z = 1.0,
       tphhl$OE1$Z = 1.0,
       tpllh$I0$Z$I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphhl$I0$Z$I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tpllh$I0$Z$I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphhl$I0$Z$I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tpllh$I1$Z$I0_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tphhl$I1$Z$I0_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tpllh$I1$Z$I0_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tphhl$I1$Z$I0_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tpllh$I2$Z$I0_EQ_0_AN_I1_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1 = 1.0,
       tphhl$I2$Z$I0_EQ_0_AN_I1_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1 = 1.0,
       tpllh$I2$Z$I0_EQ_1_AN_I1_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1 = 1.0,
       tphhl$I2$Z$I0_EQ_1_AN_I1_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1 = 1.0,
       tpllh$OE0$Z$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphhl$OE0$Z$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE1_EQ_0 = 1.0,
       tpllh$OE0$Z$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE1_EQ_0 = 1.0,
       tphhl$OE0$Z$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE1_EQ_0 = 1.0,
       tplhl$OE0$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphlh$OE0$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE1_EQ_0 = 1.0,
       tplhl$OE0$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE1_EQ_0 = 1.0,
       tphlh$OE0$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE1_EQ_0 = 1.0,
       tpllh$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_1 = 1.0,
       tphhl$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_1 = 1.0,
       tpllh$OE1$Z$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_0 = 1.0,
       tphhl$OE1$Z$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_0 = 1.0,
       tplhl$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0 = 1.0,
       tphlh$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0 = 1.0,
       tplhl$OE1$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE0_EQ_1 = 1.0,
       tphlh$OE1$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE0_EQ_1 = 1.0;

     // path delays
      (posedge OE1 => (Z +: Z)) = (1.0, 1.0);
      (negedge OE1 => (Z -: Z)) = (1.0, 1.0);

     if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && OE0 == 1'b1)
       (OE1 *> Z) = (tphlh$OE1$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE0_EQ_1, tplhl$OE1$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE0_EQ_1);
     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && OE0 == 1'b1)
       (OE1 *> Z) = (tpllh$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_1, tphhl$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_1);
     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && OE0 == 1'b0)
       (OE1 *> Z) = (tphlh$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0, tplhl$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0);
     if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && OE0 == 1'b0)
       (OE1 *> Z) = (tpllh$OE1$Z$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_0, tphhl$OE1$Z$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_0);
   //  ifnone
 //      (OE1 *> Z) = (tpllh$OE1$Z,tplhl$OE1$Z);

      (posedge OE0 => (Z +: Z)) = (1.0, 1.0);
      (negedge OE0 => (Z -: Z)) = (1.0, 1.0);
     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && OE1 == 1'b0)
       (OE0 *> Z) = (tphlh$OE0$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE1_EQ_0, tplhl$OE0$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE1_EQ_0);
     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && OE1 == 1'b0)
       (OE0 *> Z) = (tphlh$OE0$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE1_EQ_0, tplhl$OE0$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE1_EQ_0);
     if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && OE1 == 1'b0)
       (OE0 *> Z) = (tpllh$OE0$Z$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE1_EQ_0, tphhl$OE0$Z$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE1_EQ_0);
     if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && OE1 == 1'b0)
       (OE0 *> Z) = (tpllh$OE0$Z$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE1_EQ_0, tphhl$OE0$Z$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE1_EQ_0);
   //  ifnone
   //    (OE0 *> Z) = (tpllh$OE0$Z,tplhl$OE0$Z);
      (posedge I2 => (Z +: Z)) = (1.0, 1.0);
     if (I0 == 1'b1 && I1 == 1'b1 && OE0 == 1'b1 && OE1 == 1'b1)
       (I2 *> Z) = (tpllh$I2$Z$I0_EQ_1_AN_I1_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1, tphhl$I2$Z$I0_EQ_1_AN_I1_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1);
     if (I0 == 1'b0 && I1 == 1'b0 && OE0 == 1'b0 && OE1 == 1'b1)
       (I2 *> Z) = (tpllh$I2$Z$I0_EQ_0_AN_I1_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1, tphhl$I2$Z$I0_EQ_0_AN_I1_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1);
  //   ifnone
   //    (I2 *> Z) = (tpllh$I2$Z,tphhl$I2$Z);
      (posedge I1 => (Z +: Z)) = (1.0, 1.0);
     if (I0 == 1'b1 && I2 == 1'b1 && OE0 == 1'b1 && OE1 == 1'b0)
       (I1 *> Z) = (tpllh$I1$Z$I0_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0, tphhl$I1$Z$I0_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0);
     if (I0 == 1'b0 && I2 == 1'b0 && OE0 == 1'b1 && OE1 == 1'b0)
       (I1 *> Z) = (tpllh$I1$Z$I0_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0, tphhl$I1$Z$I0_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0);
  //   ifnone
  //     (I1 *> Z) = (tpllh$I1$Z,tphhl$I1$Z);
      (posedge I0 => (Z +: Z)) = (1.0, 1.0);
     if (I1 == 1'b1 && I2 == 1'b1 && OE0 == 1'b0 && OE1 == 1'b0)
       (I0 *> Z) = (tpllh$I0$Z$I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0, tphhl$I0$Z$I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0);
     if (I1 == 1'b0 && I2 == 1'b0 && OE0 == 1'b0 && OE1 == 1'b0)
       (I0 *> Z) = (tpllh$I0$Z$I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0, tphhl$I0$Z$I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0);
  //   ifnone
   //    (I0 *> Z) = (tpllh$I0$Z,tphhl$I0$Z);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_MX04D1 (Z, I0, I1, I2, I3, OE0, OE1);
input  I0 ;
input  I1 ;
input  I2 ;
input  I3 ;
input  OE0 ;
input  OE1 ;
output Z ;

   udp_mux2 (I0_out, I2, I3, OE0);
   udp_mux2 (I1_out, I0, I1, OE0);
   udp_mux2 (Z, I1_out, I0_out, OE1);

   specify
     // delay parameters
   /*  specparam
       tpllh$I0$Z = 1.0,
       tphhl$I0$Z = 1.0,
       tpllh$I1$Z = 1.0,
       tphhl$I1$Z = 1.0,
       tpllh$I2$Z = 1.0,
       tphhl$I2$Z = 1.0,
       tpllh$I3$Z = 1.0,
       tphhl$I3$Z = 1.0,
       tpllh$OE0$Z = 1.0,
       tplhl$OE0$Z = 1.0,
       tphlh$OE0$Z = 1.0,
       tphhl$OE0$Z = 1.0,
       tpllh$OE1$Z = 1.0,
       tplhl$OE1$Z = 1.0,
       tphlh$OE1$Z = 1.0,
       tphhl$OE1$Z = 1.0,
       tpllh$I0$Z$I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphhl$I0$Z$I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tpllh$I0$Z$I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphhl$I0$Z$I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tpllh$I1$Z$I0_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tphhl$I1$Z$I0_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tpllh$I1$Z$I0_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tphhl$I1$Z$I0_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tpllh$I2$Z$I0_EQ_1_AN_I1_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_1 = 1.0,
       tphhl$I2$Z$I0_EQ_1_AN_I1_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_1 = 1.0,
       tpllh$I2$Z$I0_EQ_0_AN_I1_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1 = 1.0,
       tphhl$I2$Z$I0_EQ_0_AN_I1_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1 = 1.0,
       tpllh$I3$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1 = 1.0,
       tphhl$I3$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1 = 1.0,
       tpllh$I3$Z$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_1 = 1.0,
       tphhl$I3$Z$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_1 = 1.0,
       tpllh$OE0$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_1_AN_OE1_EQ_1 = 1.0,
       tphhl$OE0$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_1_AN_OE1_EQ_1 = 1.0,
       tpllh$OE0$Z$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphhl$OE0$Z$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0 = 1.0,
       tplhl$OE0$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE1_EQ_1 = 1.0,
       tphlh$OE0$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE1_EQ_1 = 1.0,
       tplhl$OE0$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphlh$OE0$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0 = 1.0,
       tpllh$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1 = 1.0,
       tphhl$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1 = 1.0,
       tpllh$OE1$Z$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_0 = 1.0,
       tphhl$OE1$Z$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_0 = 1.0,
       tplhl$OE1$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_1 = 1.0,
       tphlh$OE1$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_1 = 1.0,
       tplhl$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0 = 1.0,
       tphlh$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0 = 1.0;

     // path delays
     if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && OE0 == 1'b1)
       (OE1 *> Z) = (tphlh$OE1$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_1, tplhl$OE1$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_1);
     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && OE0 == 1'b1)
       (OE1 *> Z) = (tpllh$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1, tphhl$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1);
     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && OE0 == 1'b0)
       (OE1 *> Z) = (tphlh$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0, tplhl$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0);
     if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && OE0 == 1'b0)
       (OE1 *> Z) = (tpllh$OE1$Z$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_0, tphhl$OE1$Z$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_0);
     ifnone
       (OE1 *> Z) = (tpllh$OE1$Z,tplhl$OE1$Z);

     if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && OE1 == 1'b1)
       (OE0 *> Z) = (tphlh$OE0$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE1_EQ_1, tplhl$OE0$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE1_EQ_1);
     if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && OE1 == 1'b1)
       (OE0 *> Z) = (tpllh$OE0$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_1_AN_OE1_EQ_1, tphhl$OE0$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_1_AN_OE1_EQ_1);
     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && OE1 == 1'b0)
       (OE0 *> Z) = (tphlh$OE0$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0, tplhl$OE0$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0);
     if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && OE1 == 1'b0)
       (OE0 *> Z) = (tpllh$OE0$Z$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0, tphhl$OE0$Z$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0);
     ifnone
       (OE0 *> Z) = (tpllh$OE0$Z,tplhl$OE0$Z);

     if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && OE0 == 1'b1 && OE1 == 1'b1)
       (I3 *> Z) = (tpllh$I3$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1, tphhl$I3$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1);
     if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && OE0 == 1'b1 && OE1 == 1'b1)
       (I3 *> Z) = (tpllh$I3$Z$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_1, tphhl$I3$Z$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_1);
     ifnone
       (I3 *> Z) = (tpllh$I3$Z,tphhl$I3$Z);

     if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b1 && OE0 == 1'b0 && OE1 == 1'b1)
       (I2 *> Z) = (tpllh$I2$Z$I0_EQ_1_AN_I1_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_1, tphhl$I2$Z$I0_EQ_1_AN_I1_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_1);
     if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b0 && OE0 == 1'b0 && OE1 == 1'b1)
       (I2 *> Z) = (tpllh$I2$Z$I0_EQ_0_AN_I1_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1, tphhl$I2$Z$I0_EQ_0_AN_I1_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1);
     ifnone
       (I2 *> Z) = (tpllh$I2$Z,tphhl$I2$Z);

     if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && OE0 == 1'b1 && OE1 == 1'b0)
       (I1 *> Z) = (tpllh$I1$Z$I0_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0, tphhl$I1$Z$I0_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0);
     if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && OE0 == 1'b1 && OE1 == 1'b0)
       (I1 *> Z) = (tpllh$I1$Z$I0_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0, tphhl$I1$Z$I0_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0);
     ifnone
       (I1 *> Z) = (tpllh$I1$Z,tphhl$I1$Z);

     if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && OE0 == 1'b0 && OE1 == 1'b0)
       (I0 *> Z) = (tpllh$I0$Z$I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0, tphhl$I0$Z$I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0);
     if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && OE0 == 1'b0 && OE1 == 1'b0)
       (I0 *> Z) = (tpllh$I0$Z$I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0, tphhl$I0$Z$I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0);
     ifnone
       (I0 *> Z) = (tpllh$I0$Z,tphhl$I0$Z);*/

   // path delays

      (posedge OE1 => (Z +: Z)) = (1.0, 1.0);
      (negedge OE1 => (Z -: Z)) = (1.0, 1.0);
      if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && OE0 == 1'b1) (OE1 +=> Z) = (1.0, 1.0);
      if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && OE0 == 1'b0) (OE1 +=> Z) = (1.0, 1.0);
      if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && OE0 == 1'b1) (OE1 -=> Z) = (1.0, 1.0);
      if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && OE0 == 1'b0) (OE1 -=> Z) = (1.0, 1.0);

      (posedge OE0 => (Z +: Z)) = (1.0, 1.0);
      (negedge OE0 => (Z -: Z)) = (1.0, 1.0);
      if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && OE1 == 1'b0) (OE0 +=> Z) = (1.0, 1.0);
      if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && OE1 == 1'b1) (OE0 +=> Z) = (1.0, 1.0);
      if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && OE1 == 1'b0) (OE0 -=> Z) = (1.0, 1.0);
      if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && OE1 == 1'b1) (OE0 -=> Z) = (1.0, 1.0);

      (posedge I3 => (Z +: Z)) = (1.0, 1.0);
      //(negedge I3 => (Z -: Z)) = (1.0, 1.0);
      if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && OE0 == 1'b1 && OE1 == 1'b1) (I3 +=> Z) = (1.0, 1.0);
      if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && OE0 == 1'b1 && OE1 == 1'b1) (I3 +=> Z) = (1.0, 1.0);

      (posedge I2 => (Z +: Z)) = (1.0, 1.0);
      if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b1 && OE0 == 1'b0 && OE1 == 1'b1) (I2 +=> Z) = (1.0, 1.0);
      if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b0 && OE0 == 1'b0 && OE1 == 1'b1) (I2 +=> Z) = (1.0, 1.0);

      (posedge I1 => (Z +: Z)) = (1.0, 1.0);
      if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && OE0 == 1'b1 && OE1 == 1'b0) (I1 +=> Z) = (1.0, 1.0);
      if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && OE0 == 1'b1 && OE1 == 1'b0) (I1 +=> Z) = (1.0, 1.0);

      (posedge I0 => (Z +: Z)) = (1.0, 1.0);
      if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && OE0 == 1'b0 && OE1 == 1'b0) (I0 +=> Z) = (1.0, 1.0);
      if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && OE0 == 1'b0 && OE1 == 1'b0) (I0 +=> Z) = (1.0, 1.0);



   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_MX04D2 (Z, I0, I1, I2, I3, OE0, OE1);
input  I0 ;
input  I1 ;
input  I2 ;
input  I3 ;
input  OE0 ;
input  OE1 ;
output Z ;

   udp_mux2 (I0_out, I2, I3, OE0);
   udp_mux2 (I1_out, I0, I1, OE0);
   udp_mux2 (Z, I1_out, I0_out, OE1);

   specify
     // delay parameters
 /*    specparam
       tpllh$I0$Z = 1.0,
       tphhl$I0$Z = 1.0,
       tpllh$I1$Z = 1.0,
       tphhl$I1$Z = 1.0,
       tpllh$I2$Z = 1.0,
       tphhl$I2$Z = 1.0,
       tpllh$I3$Z = 1.0,
       tphhl$I3$Z = 1.0,
       tpllh$OE0$Z = 1.0,
       tplhl$OE0$Z = 1.0,
       tphlh$OE0$Z = 1.0,
       tphhl$OE0$Z = 1.0,
       tpllh$OE1$Z = 1.0,
       tplhl$OE1$Z = 1.0,
       tphlh$OE1$Z = 1.0,
       tphhl$OE1$Z = 1.0,
       tpllh$I0$Z$I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphhl$I0$Z$I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tpllh$I0$Z$I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphhl$I0$Z$I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tpllh$I1$Z$I0_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tphhl$I1$Z$I0_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tpllh$I1$Z$I0_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tphhl$I1$Z$I0_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tpllh$I2$Z$I0_EQ_1_AN_I1_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_1 = 1.0,
       tphhl$I2$Z$I0_EQ_1_AN_I1_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_1 = 1.0,
       tpllh$I2$Z$I0_EQ_0_AN_I1_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1 = 1.0,
       tphhl$I2$Z$I0_EQ_0_AN_I1_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1 = 1.0,
       tpllh$I3$Z$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_1 = 1.0,
       tphhl$I3$Z$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_1 = 1.0,
       tpllh$I3$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1 = 1.0,
       tphhl$I3$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1 = 1.0,
       tpllh$OE0$Z$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphhl$OE0$Z$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0 = 1.0,
       tpllh$OE0$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_1_AN_OE1_EQ_1 = 1.0,
       tphhl$OE0$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_1_AN_OE1_EQ_1 = 1.0,
       tplhl$OE0$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphlh$OE0$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0 = 1.0,
       tplhl$OE0$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE1_EQ_1 = 1.0,
       tphlh$OE0$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE1_EQ_1 = 1.0,
       tpllh$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1 = 1.0,
       tphhl$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1 = 1.0,
       tpllh$OE1$Z$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_0 = 1.0,
       tphhl$OE1$Z$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_0 = 1.0,
       tplhl$OE1$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_1 = 1.0,
       tphlh$OE1$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_1 = 1.0,
       tplhl$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0 = 1.0,
       tphlh$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0 = 1.0;

     // path delays
     if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && OE0 == 1'b1)
       (OE1 *> Z) = (tphlh$OE1$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_1, tplhl$OE1$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_1);
     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && OE0 == 1'b1)
       (OE1 *> Z) = (tpllh$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1, tphhl$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1);
     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && OE0 == 1'b0)
       (OE1 *> Z) = (tphlh$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0, tplhl$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0);
     if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && OE0 == 1'b0)
       (OE1 *> Z) = (tpllh$OE1$Z$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_0, tphhl$OE1$Z$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_0);
     ifnone
       (OE1 *> Z) = (tpllh$OE1$Z,tplhl$OE1$Z);

     if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && OE1 == 1'b1)
       (OE0 *> Z) = (tphlh$OE0$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE1_EQ_1, tplhl$OE0$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE1_EQ_1);
     if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && OE1 == 1'b1)
       (OE0 *> Z) = (tpllh$OE0$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_1_AN_OE1_EQ_1, tphhl$OE0$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_1_AN_OE1_EQ_1);
     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && OE1 == 1'b0)
       (OE0 *> Z) = (tphlh$OE0$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0, tplhl$OE0$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0);
     if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && OE1 == 1'b0)
       (OE0 *> Z) = (tpllh$OE0$Z$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0, tphhl$OE0$Z$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0);
     ifnone
       (OE0 *> Z) = (tpllh$OE0$Z,tplhl$OE0$Z);

     if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && OE0 == 1'b1 && OE1 == 1'b1)
       (I3 *> Z) = (tpllh$I3$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1, tphhl$I3$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1);
     if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && OE0 == 1'b1 && OE1 == 1'b1)
       (I3 *> Z) = (tpllh$I3$Z$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_1, tphhl$I3$Z$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_1);
     ifnone
       (I3 *> Z) = (tpllh$I3$Z,tphhl$I3$Z);

     if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b1 && OE0 == 1'b0 && OE1 == 1'b1)
       (I2 *> Z) = (tpllh$I2$Z$I0_EQ_1_AN_I1_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_1, tphhl$I2$Z$I0_EQ_1_AN_I1_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_1);
     if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b0 && OE0 == 1'b0 && OE1 == 1'b1)
       (I2 *> Z) = (tpllh$I2$Z$I0_EQ_0_AN_I1_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1, tphhl$I2$Z$I0_EQ_0_AN_I1_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1);
     ifnone
       (I2 *> Z) = (tpllh$I2$Z,tphhl$I2$Z);

     if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && OE0 == 1'b1 && OE1 == 1'b0)
       (I1 *> Z) = (tpllh$I1$Z$I0_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0, tphhl$I1$Z$I0_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0);
     if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && OE0 == 1'b1 && OE1 == 1'b0)
       (I1 *> Z) = (tpllh$I1$Z$I0_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0, tphhl$I1$Z$I0_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0);
     ifnone
       (I1 *> Z) = (tpllh$I1$Z,tphhl$I1$Z);

     if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && OE0 == 1'b0 && OE1 == 1'b0)
       (I0 *> Z) = (tpllh$I0$Z$I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0, tphhl$I0$Z$I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0);
     if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && OE0 == 1'b0 && OE1 == 1'b0)
       (I0 *> Z) = (tpllh$I0$Z$I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0, tphhl$I0$Z$I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0);
     ifnone
       (I0 *> Z) = (tpllh$I0$Z,tphhl$I0$Z);*/

   // path delays

      (posedge OE1 => (Z +: Z)) = (1.0, 1.0);
      (negedge OE1 => (Z -: Z)) = (1.0, 1.0);
      if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && OE0 == 1'b1) (OE1 +=> Z) = (1.0, 1.0);
      if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && OE0 == 1'b0) (OE1 +=> Z) = (1.0, 1.0);
      if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && OE0 == 1'b1) (OE1 -=> Z) = (1.0, 1.0);
      if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && OE0 == 1'b0) (OE1 -=> Z) = (1.0, 1.0);

      (posedge OE0 => (Z +: Z)) = (1.0, 1.0);
      (negedge OE0 => (Z -: Z)) = (1.0, 1.0);
      if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && OE1 == 1'b0) (OE0 +=> Z) = (1.0, 1.0);
      if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && OE1 == 1'b1) (OE0 +=> Z) = (1.0, 1.0);
      if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && OE1 == 1'b0) (OE0 -=> Z) = (1.0, 1.0);
      if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && OE1 == 1'b1) (OE0 -=> Z) = (1.0, 1.0);

      (posedge I3 => (Z +: Z)) = (1.0, 1.0);
      //(negedge I3 => (Z -: Z)) = (1.0, 1.0);
      if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && OE0 == 1'b1 && OE1 == 1'b1) (I3 +=> Z) = (1.0, 1.0);
      if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && OE0 == 1'b1 && OE1 == 1'b1) (I3 +=> Z) = (1.0, 1.0);

      (posedge I2 => (Z +: Z)) = (1.0, 1.0);
      if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b1 && OE0 == 1'b0 && OE1 == 1'b1) (I2 +=> Z) = (1.0, 1.0);
      if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b0 && OE0 == 1'b0 && OE1 == 1'b1) (I2 +=> Z) = (1.0, 1.0);

      (posedge I1 => (Z +: Z)) = (1.0, 1.0);
      if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && OE0 == 1'b1 && OE1 == 1'b0) (I1 +=> Z) = (1.0, 1.0);
      if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && OE0 == 1'b1 && OE1 == 1'b0) (I1 +=> Z) = (1.0, 1.0);

      (posedge I0 => (Z +: Z)) = (1.0, 1.0);
      if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && OE0 == 1'b0 && OE1 == 1'b0) (I0 +=> Z) = (1.0, 1.0);
      if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && OE0 == 1'b0 && OE1 == 1'b0) (I0 +=> Z) = (1.0, 1.0);





   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_MX04D4 (Z, I0, I1, I2, I3, OE0, OE1);
input  I0 ;
input  I1 ;
input  I2 ;
input  I3 ;
input  OE0 ;
input  OE1 ;
output Z ;

   udp_mux2 (I0_out, I2, I3, OE0);
   udp_mux2 (I1_out, I0, I1, OE0);
   udp_mux2 (Z, I1_out, I0_out, OE1);

   specify
     // delay parameters
/*     specparam
       tpllh$I0$Z = 1.0,
       tphhl$I0$Z = 1.0,
       tpllh$I1$Z = 1.0,
       tphhl$I1$Z = 1.0,
       tpllh$I2$Z = 1.0,
       tphhl$I2$Z = 1.0,
       tpllh$I3$Z = 1.0,
       tphhl$I3$Z = 1.0,
       tpllh$OE0$Z = 1.0,
       tplhl$OE0$Z = 1.0,
       tphlh$OE0$Z = 1.0,
       tphhl$OE0$Z = 1.0,
       tpllh$OE1$Z = 1.0,
       tplhl$OE1$Z = 1.0,
       tphlh$OE1$Z = 1.0,
       tphhl$OE1$Z = 1.0,
       tpllh$I0$Z$I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphhl$I0$Z$I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tpllh$I0$Z$I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphhl$I0$Z$I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tpllh$I1$Z$I0_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tphhl$I1$Z$I0_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tpllh$I1$Z$I0_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tphhl$I1$Z$I0_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tpllh$I2$Z$I0_EQ_1_AN_I1_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_1 = 1.0,
       tphhl$I2$Z$I0_EQ_1_AN_I1_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_1 = 1.0,
       tpllh$I2$Z$I0_EQ_0_AN_I1_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1 = 1.0,
       tphhl$I2$Z$I0_EQ_0_AN_I1_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1 = 1.0,
       tpllh$I3$Z$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_1 = 1.0,
       tphhl$I3$Z$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_1 = 1.0,
       tpllh$I3$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1 = 1.0,
       tphhl$I3$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1 = 1.0,
       tpllh$OE0$Z$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphhl$OE0$Z$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0 = 1.0,
       tpllh$OE0$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_1_AN_OE1_EQ_1 = 1.0,
       tphhl$OE0$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_1_AN_OE1_EQ_1 = 1.0,
       tplhl$OE0$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphlh$OE0$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0 = 1.0,
       tplhl$OE0$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE1_EQ_1 = 1.0,
       tphlh$OE0$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE1_EQ_1 = 1.0,
       tpllh$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1 = 1.0,
       tphhl$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1 = 1.0,
       tpllh$OE1$Z$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_0 = 1.0,
       tphhl$OE1$Z$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_0 = 1.0,
       tplhl$OE1$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_1 = 1.0,
       tphlh$OE1$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_1 = 1.0,
       tplhl$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0 = 1.0,
       tphlh$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0 = 1.0;

     // path delays
     if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && OE0 == 1'b1)
       (OE1 *> Z) = (tphlh$OE1$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_1, tplhl$OE1$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_1);
     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && OE0 == 1'b1)
       (OE1 *> Z) = (tpllh$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1, tphhl$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1);
     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && OE0 == 1'b0)
       (OE1 *> Z) = (tphlh$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0, tplhl$OE1$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0);
     if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && OE0 == 1'b0)
       (OE1 *> Z) = (tpllh$OE1$Z$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_0, tphhl$OE1$Z$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_0);
     ifnone
       (OE1 *> Z) = (tpllh$OE1$Z,tplhl$OE1$Z);

     if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && OE1 == 1'b1)
       (OE0 *> Z) = (tphlh$OE0$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE1_EQ_1, tplhl$OE0$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE1_EQ_1);
     if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && OE1 == 1'b1)
       (OE0 *> Z) = (tpllh$OE0$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_1_AN_OE1_EQ_1, tphhl$OE0$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_1_AN_OE1_EQ_1);
     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && OE1 == 1'b0)
       (OE0 *> Z) = (tphlh$OE0$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0, tplhl$OE0$Z$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0);
     if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && OE1 == 1'b0)
       (OE0 *> Z) = (tpllh$OE0$Z$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0, tphhl$OE0$Z$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0);
     ifnone
       (OE0 *> Z) = (tpllh$OE0$Z,tplhl$OE0$Z);

     if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && OE0 == 1'b1 && OE1 == 1'b1)
       (I3 *> Z) = (tpllh$I3$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1, tphhl$I3$Z$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1);
     if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && OE0 == 1'b1 && OE1 == 1'b1)
       (I3 *> Z) = (tpllh$I3$Z$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_1, tphhl$I3$Z$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_1);
     ifnone
       (I3 *> Z) = (tpllh$I3$Z,tphhl$I3$Z);

     if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b1 && OE0 == 1'b0 && OE1 == 1'b1)
       (I2 *> Z) = (tpllh$I2$Z$I0_EQ_1_AN_I1_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_1, tphhl$I2$Z$I0_EQ_1_AN_I1_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_1);
     if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b0 && OE0 == 1'b0 && OE1 == 1'b1)
       (I2 *> Z) = (tpllh$I2$Z$I0_EQ_0_AN_I1_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1, tphhl$I2$Z$I0_EQ_0_AN_I1_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1);
     ifnone
       (I2 *> Z) = (tpllh$I2$Z,tphhl$I2$Z);

     if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && OE0 == 1'b1 && OE1 == 1'b0)
       (I1 *> Z) = (tpllh$I1$Z$I0_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0, tphhl$I1$Z$I0_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0);
     if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && OE0 == 1'b1 && OE1 == 1'b0)
       (I1 *> Z) = (tpllh$I1$Z$I0_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0, tphhl$I1$Z$I0_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0);
     ifnone
       (I1 *> Z) = (tpllh$I1$Z,tphhl$I1$Z);

     if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && OE0 == 1'b0 && OE1 == 1'b0)
       (I0 *> Z) = (tpllh$I0$Z$I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0, tphhl$I0$Z$I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0);
     if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && OE0 == 1'b0 && OE1 == 1'b0)
       (I0 *> Z) = (tpllh$I0$Z$I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0, tphhl$I0$Z$I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0);
     ifnone
       (I0 *> Z) = (tpllh$I0$Z,tphhl$I0$Z);*/

   // path delays

      (posedge OE1 => (Z +: Z)) = (1.0, 1.0);
      (negedge OE1 => (Z -: Z)) = (1.0, 1.0);
      if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && OE0 == 1'b1) (OE1 +=> Z) = (1.0, 1.0);
      if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && OE0 == 1'b0) (OE1 +=> Z) = (1.0, 1.0);
      if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && OE0 == 1'b1) (OE1 -=> Z) = (1.0, 1.0);
      if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && OE0 == 1'b0) (OE1 -=> Z) = (1.0, 1.0);

      (posedge OE0 => (Z +: Z)) = (1.0, 1.0);
      (negedge OE0 => (Z -: Z)) = (1.0, 1.0);
      if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && OE1 == 1'b0) (OE0 +=> Z) = (1.0, 1.0);
      if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && OE1 == 1'b1) (OE0 +=> Z) = (1.0, 1.0);
      if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && OE1 == 1'b0) (OE0 -=> Z) = (1.0, 1.0);
      if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && OE1 == 1'b1) (OE0 -=> Z) = (1.0, 1.0);

      (posedge I3 => (Z +: Z)) = (1.0, 1.0);
      //(negedge I3 => (Z -: Z)) = (1.0, 1.0);
      if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && OE0 == 1'b1 && OE1 == 1'b1) (I3 +=> Z) = (1.0, 1.0);
      if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && OE0 == 1'b1 && OE1 == 1'b1) (I3 +=> Z) = (1.0, 1.0);

      (posedge I2 => (Z +: Z)) = (1.0, 1.0);
      if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b1 && OE0 == 1'b0 && OE1 == 1'b1) (I2 +=> Z) = (1.0, 1.0);
      if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b0 && OE0 == 1'b0 && OE1 == 1'b1) (I2 +=> Z) = (1.0, 1.0);

      (posedge I1 => (Z +: Z)) = (1.0, 1.0);
      if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && OE0 == 1'b1 && OE1 == 1'b0) (I1 +=> Z) = (1.0, 1.0);
      if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && OE0 == 1'b1 && OE1 == 1'b0) (I1 +=> Z) = (1.0, 1.0);

      (posedge I0 => (Z +: Z)) = (1.0, 1.0);
      if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && OE0 == 1'b0 && OE1 == 1'b0) (I0 +=> Z) = (1.0, 1.0);
      if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && OE0 == 1'b0 && OE1 == 1'b0) (I0 +=> Z) = (1.0, 1.0);



   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_MXI2D1 (ZN, I0, I1, OE);
input  I0 ;
input  I1 ;
input  OE ;
output ZN ;

   udp_mux2 (I0_out, I0, I1, OE);
   not (ZN, I0_out);

   specify
     // delay parameters
     specparam
       tplhl$I0$ZN = 1.0,
       tphlh$I0$ZN = 1.0,
       tplhl$I1$ZN = 1.0,
       tphlh$I1$ZN = 1.0,
       tpllh$OE$ZN = 1.0,
       tplhl$OE$ZN = 1.0,
       tphlh$OE$ZN = 1.0,
       tphhl$OE$ZN = 1.0,
       tplhl$I0$ZN$I1_EQ_1_AN_OE_EQ_0 = 1.0,
       tphlh$I0$ZN$I1_EQ_1_AN_OE_EQ_0 = 1.0,
       tplhl$I0$ZN$I1_EQ_0_AN_OE_EQ_0 = 1.0,
       tphlh$I0$ZN$I1_EQ_0_AN_OE_EQ_0 = 1.0,
       tplhl$I1$ZN$I0_EQ_0_AN_OE_EQ_1 = 1.0,
       tphlh$I1$ZN$I0_EQ_0_AN_OE_EQ_1 = 1.0,
       tplhl$I1$ZN$I0_EQ_1_AN_OE_EQ_1 = 1.0,
       tphlh$I1$ZN$I0_EQ_1_AN_OE_EQ_1 = 1.0;

     // path delays
     (posedge OE *> (ZN +: !I1)) = (tpllh$OE$ZN, tplhl$OE$ZN);
     (negedge OE *> (ZN +: !I0)) = (tphlh$OE$ZN, tphhl$OE$ZN);
     if (I0 == 1'b1 && OE == 1'b1)
       (I1 *> ZN) = (tphlh$I1$ZN$I0_EQ_1_AN_OE_EQ_1, tplhl$I1$ZN$I0_EQ_1_AN_OE_EQ_1);
     if (I0 == 1'b0 && OE == 1'b1)
       (I1 *> ZN) = (tphlh$I1$ZN$I0_EQ_0_AN_OE_EQ_1, tplhl$I1$ZN$I0_EQ_0_AN_OE_EQ_1);
     ifnone
       (I1 *> ZN) = (tphlh$I1$ZN,tplhl$I1$ZN);

     if (I1 == 1'b1 && OE == 1'b0)
       (I0 *> ZN) = (tphlh$I0$ZN$I1_EQ_1_AN_OE_EQ_0, tplhl$I0$ZN$I1_EQ_1_AN_OE_EQ_0);
     if (I1 == 1'b0 && OE == 1'b0)
       (I0 *> ZN) = (tphlh$I0$ZN$I1_EQ_0_AN_OE_EQ_0, tplhl$I0$ZN$I1_EQ_0_AN_OE_EQ_0);
     ifnone
       (I0 *> ZN) = (tphlh$I0$ZN,tplhl$I0$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_MXI2D2 (ZN, I0, I1, OE);
input  I0 ;
input  I1 ;
input  OE ;
output ZN ;

   udp_mux2 (I0_out, I0, I1, OE);
   not (ZN, I0_out);

   specify
     // delay parameters
     specparam
       tplhl$I0$ZN = 1.0,
       tphlh$I0$ZN = 1.0,
       tplhl$I1$ZN = 1.0,
       tphlh$I1$ZN = 1.0,
       tpllh$OE$ZN = 1.0,
       tplhl$OE$ZN = 1.0,
       tphlh$OE$ZN = 1.0,
       tphhl$OE$ZN = 1.0,
       tplhl$I0$ZN$I1_EQ_1_AN_OE_EQ_0 = 1.0,
       tphlh$I0$ZN$I1_EQ_1_AN_OE_EQ_0 = 1.0,
       tplhl$I0$ZN$I1_EQ_0_AN_OE_EQ_0 = 1.0,
       tphlh$I0$ZN$I1_EQ_0_AN_OE_EQ_0 = 1.0,
       tplhl$I1$ZN$I0_EQ_1_AN_OE_EQ_1 = 1.0,
       tphlh$I1$ZN$I0_EQ_1_AN_OE_EQ_1 = 1.0,
       tplhl$I1$ZN$I0_EQ_0_AN_OE_EQ_1 = 1.0,
       tphlh$I1$ZN$I0_EQ_0_AN_OE_EQ_1 = 1.0;

     // path delays
     (posedge OE *> (ZN +: !I1)) = (tpllh$OE$ZN, tplhl$OE$ZN);
     (negedge OE *> (ZN +: !I0)) = (tphlh$OE$ZN, tphhl$OE$ZN);
     if (I0 == 1'b1 && OE == 1'b1)
       (I1 *> ZN) = (tphlh$I1$ZN$I0_EQ_1_AN_OE_EQ_1, tplhl$I1$ZN$I0_EQ_1_AN_OE_EQ_1);
     if (I0 == 1'b0 && OE == 1'b1)
       (I1 *> ZN) = (tphlh$I1$ZN$I0_EQ_0_AN_OE_EQ_1, tplhl$I1$ZN$I0_EQ_0_AN_OE_EQ_1);
     ifnone
       (I1 *> ZN) = (tphlh$I1$ZN,tplhl$I1$ZN);

     if (I1 == 1'b1 && OE == 1'b0)
       (I0 *> ZN) = (tphlh$I0$ZN$I1_EQ_1_AN_OE_EQ_0, tplhl$I0$ZN$I1_EQ_1_AN_OE_EQ_0);
     if (I1 == 1'b0 && OE == 1'b0)
       (I0 *> ZN) = (tphlh$I0$ZN$I1_EQ_0_AN_OE_EQ_0, tplhl$I0$ZN$I1_EQ_0_AN_OE_EQ_0);
     ifnone
       (I0 *> ZN) = (tphlh$I0$ZN,tplhl$I0$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_MXI2D4 (ZN, I0, I1, OE);
input  I0 ;
input  I1 ;
input  OE ;
output ZN ;

   udp_mux2 (I0_out, I0, I1, OE);
   not (ZN, I0_out);

   specify
     // delay parameters
     specparam
       tplhl$I0$ZN = 1.0,
       tphlh$I0$ZN = 1.0,
       tplhl$I1$ZN = 1.0,
       tphlh$I1$ZN = 1.0,
       tpllh$OE$ZN = 1.0,
       tplhl$OE$ZN = 1.0,
       tphlh$OE$ZN = 1.0,
       tphhl$OE$ZN = 1.0,
       tplhl$I0$ZN$I1_EQ_1_AN_OE_EQ_0 = 1.0,
       tphlh$I0$ZN$I1_EQ_1_AN_OE_EQ_0 = 1.0,
       tplhl$I0$ZN$I1_EQ_0_AN_OE_EQ_0 = 1.0,
       tphlh$I0$ZN$I1_EQ_0_AN_OE_EQ_0 = 1.0,
       tplhl$I1$ZN$I0_EQ_0_AN_OE_EQ_1 = 1.0,
       tphlh$I1$ZN$I0_EQ_0_AN_OE_EQ_1 = 1.0,
       tplhl$I1$ZN$I0_EQ_1_AN_OE_EQ_1 = 1.0,
       tphlh$I1$ZN$I0_EQ_1_AN_OE_EQ_1 = 1.0;

     // path delays
     (posedge OE *> (ZN +: !I1)) = (tpllh$OE$ZN, tplhl$OE$ZN);
     (negedge OE *> (ZN +: !I0)) = (tphlh$OE$ZN, tphhl$OE$ZN);
     if (I0 == 1'b1 && OE == 1'b1)
       (I1 *> ZN) = (tphlh$I1$ZN$I0_EQ_1_AN_OE_EQ_1, tplhl$I1$ZN$I0_EQ_1_AN_OE_EQ_1);
     if (I0 == 1'b0 && OE == 1'b1)
       (I1 *> ZN) = (tphlh$I1$ZN$I0_EQ_0_AN_OE_EQ_1, tplhl$I1$ZN$I0_EQ_0_AN_OE_EQ_1);
     ifnone
       (I1 *> ZN) = (tphlh$I1$ZN,tplhl$I1$ZN);

     if (I1 == 1'b1 && OE == 1'b0)
       (I0 *> ZN) = (tphlh$I0$ZN$I1_EQ_1_AN_OE_EQ_0, tplhl$I0$ZN$I1_EQ_1_AN_OE_EQ_0);
     if (I1 == 1'b0 && OE == 1'b0)
       (I0 *> ZN) = (tphlh$I0$ZN$I1_EQ_0_AN_OE_EQ_0, tplhl$I0$ZN$I1_EQ_0_AN_OE_EQ_0);
     ifnone
       (I0 *> ZN) = (tphlh$I0$ZN,tplhl$I0$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_MXI3D1 (ZN, I0, I1, I2, OE0, OE1);
input  I0 ;
input  I1 ;
input  I2 ;
input  OE0 ;
input  OE1 ;
output ZN ;

   udp_mux2 (I0_out, I0, I1, OE0);
   udp_mux2 (I1_out, I0_out, I2, OE1);
   not (ZN, I1_out);

   specify
     // delay parameters
     specparam
       tplhl$I0$ZN = 1.0,
       tphlh$I0$ZN = 1.0,
       tplhl$I1$ZN = 1.0,
       tphlh$I1$ZN = 1.0,
       tplhl$I2$ZN = 1.0,
       tphlh$I2$ZN = 1.0,
       tpllh$OE0$ZN = 1.0,
       tplhl$OE0$ZN = 1.0,
       tphlh$OE0$ZN = 1.0,
       tphhl$OE0$ZN = 1.0,
       tpllh$OE1$ZN = 1.0,
       tplhl$OE1$ZN = 1.0,
       tphlh$OE1$ZN = 1.0,
       tphhl$OE1$ZN = 1.0,
       tplhl$I0$ZN$I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphlh$I0$ZN$I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tplhl$I0$ZN$I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphlh$I0$ZN$I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tplhl$I1$ZN$I0_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tphlh$I1$ZN$I0_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tplhl$I1$ZN$I0_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tphlh$I1$ZN$I0_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tplhl$I2$ZN$I0_EQ_0_AN_I1_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1 = 1.0,
       tphlh$I2$ZN$I0_EQ_0_AN_I1_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1 = 1.0,
       tplhl$I2$ZN$I0_EQ_1_AN_I1_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1 = 1.0,
       tphlh$I2$ZN$I0_EQ_1_AN_I1_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1 = 1.0,
       tpllh$OE0$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphhl$OE0$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE1_EQ_0 = 1.0,
       tpllh$OE0$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE1_EQ_0 = 1.0,
       tphhl$OE0$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE1_EQ_0 = 1.0,
       tplhl$OE0$ZN$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphlh$OE0$ZN$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE1_EQ_0 = 1.0,
       tplhl$OE0$ZN$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE1_EQ_0 = 1.0,
       tphlh$OE0$ZN$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE1_EQ_0 = 1.0,
       tpllh$OE1$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE0_EQ_1 = 1.0,
       tphhl$OE1$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE0_EQ_1 = 1.0,
       tpllh$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0 = 1.0,
       tphhl$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0 = 1.0,
       tplhl$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_1 = 1.0,
       tphlh$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_1 = 1.0,
       tplhl$OE1$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_0 = 1.0,
       tphlh$OE1$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_0 = 1.0;

     // path delays

      (posedge OE1 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge OE1 => (ZN -: ZN)) = (1.0, 1.0);

     if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && OE0 == 1'b1)
       (OE1 *> ZN) = (tpllh$OE1$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE0_EQ_1, tphhl$OE1$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE0_EQ_1);
     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && OE0 == 1'b1)
       (OE1 *> ZN) = (tphlh$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_1, tplhl$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_1);
     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && OE0 == 1'b0)
       (OE1 *> ZN) = (tpllh$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0, tphhl$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0);
     if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && OE0 == 1'b0)
       (OE1 *> ZN) = (tphlh$OE1$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_0, tplhl$OE1$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_0);
    // ifnone
    //   (OE1 *> ZN) = (tpllh$OE1$ZN,tplhl$OE1$ZN);
    
      (posedge OE0 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge OE0 => (ZN -: ZN)) = (1.0, 1.0);


     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && OE1 == 1'b0)
       (OE0 *> ZN) = (tpllh$OE0$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE1_EQ_0, tphhl$OE0$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE1_EQ_0);
     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && OE1 == 1'b0)
       (OE0 *> ZN) = (tpllh$OE0$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE1_EQ_0, tphhl$OE0$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE1_EQ_0);
     if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && OE1 == 1'b0)
       (OE0 *> ZN) = (tphlh$OE0$ZN$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE1_EQ_0, tplhl$OE0$ZN$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE1_EQ_0);
     if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && OE1 == 1'b0)
       (OE0 *> ZN) = (tphlh$OE0$ZN$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE1_EQ_0, tplhl$OE0$ZN$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE1_EQ_0);
   //  ifnone
    //   (OE0 *> ZN) = (tpllh$OE0$ZN,tplhl$OE0$ZN);

(negedge I2 => (ZN -: ZN)) = (1.0, 1.0);
     if (I0 == 1'b1 && I1 == 1'b1 && OE0 == 1'b1 && OE1 == 1'b1)
       (I2 *> ZN) = (tphlh$I2$ZN$I0_EQ_1_AN_I1_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1, tplhl$I2$ZN$I0_EQ_1_AN_I1_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1);
     if (I0 == 1'b0 && I1 == 1'b0 && OE0 == 1'b0 && OE1 == 1'b1)
       (I2 *> ZN) = (tphlh$I2$ZN$I0_EQ_0_AN_I1_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1, tplhl$I2$ZN$I0_EQ_0_AN_I1_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1);
  //   ifnone
 //      (I2 *> ZN) = (tphlh$I2$ZN,tplhl$I2$ZN);

(negedge I1 => (ZN -: ZN)) = (1.0, 1.0);
     if (I0 == 1'b1 && I2 == 1'b1 && OE0 == 1'b1 && OE1 == 1'b0)
       (I1 *> ZN) = (tphlh$I1$ZN$I0_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0, tplhl$I1$ZN$I0_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0);
     if (I0 == 1'b0 && I2 == 1'b0 && OE0 == 1'b1 && OE1 == 1'b0)
       (I1 *> ZN) = (tphlh$I1$ZN$I0_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0, tplhl$I1$ZN$I0_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0);
 //    ifnone
   //    (I1 *> ZN) = (tphlh$I1$ZN,tplhl$I1$ZN);
(negedge I0 => (ZN -: ZN)) = (1.0, 1.0);
     if (I1 == 1'b1 && I2 == 1'b1 && OE0 == 1'b0 && OE1 == 1'b0)
       (I0 *> ZN) = (tphlh$I0$ZN$I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0, tplhl$I0$ZN$I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0);
     if (I1 == 1'b0 && I2 == 1'b0 && OE0 == 1'b0 && OE1 == 1'b0)
       (I0 *> ZN) = (tphlh$I0$ZN$I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0, tplhl$I0$ZN$I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0);
    // ifnone
  //     (I0 *> ZN) = (tphlh$I0$ZN,tplhl$I0$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_MXI3D2 (ZN, I0, I1, I2, OE0, OE1);
input  I0 ;
input  I1 ;
input  I2 ;
input  OE0 ;
input  OE1 ;
output ZN ;

   udp_mux2 (I0_out, I0, I1, OE0);
   udp_mux2 (I1_out, I0_out, I2, OE1);
   not (ZN, I1_out);

   specify
     // delay parameters
     specparam
       tplhl$I0$ZN = 1.0,
       tphlh$I0$ZN = 1.0,
       tplhl$I1$ZN = 1.0,
       tphlh$I1$ZN = 1.0,
       tplhl$I2$ZN = 1.0,
       tphlh$I2$ZN = 1.0,
       tpllh$OE0$ZN = 1.0,
       tplhl$OE0$ZN = 1.0,
       tphlh$OE0$ZN = 1.0,
       tphhl$OE0$ZN = 1.0,
       tpllh$OE1$ZN = 1.0,
       tplhl$OE1$ZN = 1.0,
       tphlh$OE1$ZN = 1.0,
       tphhl$OE1$ZN = 1.0,
       tplhl$I0$ZN$I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphlh$I0$ZN$I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tplhl$I0$ZN$I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphlh$I0$ZN$I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tplhl$I1$ZN$I0_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tphlh$I1$ZN$I0_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tplhl$I1$ZN$I0_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tphlh$I1$ZN$I0_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tplhl$I2$ZN$I0_EQ_1_AN_I1_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1 = 1.0,
       tphlh$I2$ZN$I0_EQ_1_AN_I1_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1 = 1.0,
       tplhl$I2$ZN$I0_EQ_0_AN_I1_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1 = 1.0,
       tphlh$I2$ZN$I0_EQ_0_AN_I1_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1 = 1.0,
       tpllh$OE0$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphhl$OE0$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE1_EQ_0 = 1.0,
       tpllh$OE0$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE1_EQ_0 = 1.0,
       tphhl$OE0$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE1_EQ_0 = 1.0,
       tplhl$OE0$ZN$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphlh$OE0$ZN$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE1_EQ_0 = 1.0,
       tplhl$OE0$ZN$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE1_EQ_0 = 1.0,
       tphlh$OE0$ZN$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE1_EQ_0 = 1.0,
       tpllh$OE1$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE0_EQ_1 = 1.0,
       tphhl$OE1$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE0_EQ_1 = 1.0,
       tpllh$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0 = 1.0,
       tphhl$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0 = 1.0,
       tplhl$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_1 = 1.0,
       tphlh$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_1 = 1.0,
       tplhl$OE1$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_0 = 1.0,
       tphlh$OE1$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_0 = 1.0;

     // path delays
      (posedge OE1 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge OE1 => (ZN -: ZN)) = (1.0, 1.0);

     if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && OE0 == 1'b1)
       (OE1 *> ZN) = (tpllh$OE1$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE0_EQ_1, tphhl$OE1$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE0_EQ_1);
     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && OE0 == 1'b1)
       (OE1 *> ZN) = (tphlh$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_1, tplhl$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_1);
     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && OE0 == 1'b0)
       (OE1 *> ZN) = (tpllh$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0, tphhl$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0);
     if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && OE0 == 1'b0)
       (OE1 *> ZN) = (tphlh$OE1$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_0, tplhl$OE1$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_0);
   //  ifnone
   //    (OE1 *> ZN) = (tpllh$OE1$ZN,tplhl$OE1$ZN);
      (posedge OE0 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge OE0 => (ZN -: ZN)) = (1.0, 1.0);

     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && OE1 == 1'b0)
       (OE0 *> ZN) = (tpllh$OE0$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE1_EQ_0, tphhl$OE0$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE1_EQ_0);
     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && OE1 == 1'b0)
       (OE0 *> ZN) = (tpllh$OE0$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE1_EQ_0, tphhl$OE0$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE1_EQ_0);
     if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && OE1 == 1'b0)
       (OE0 *> ZN) = (tphlh$OE0$ZN$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE1_EQ_0, tplhl$OE0$ZN$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE1_EQ_0);
     if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && OE1 == 1'b0)
       (OE0 *> ZN) = (tphlh$OE0$ZN$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE1_EQ_0, tplhl$OE0$ZN$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE1_EQ_0);
  //   ifnone
    //   (OE0 *> ZN) = (tpllh$OE0$ZN,tplhl$OE0$ZN);
(negedge I2 => (ZN -: ZN)) = (1.0, 1.0);
     if (I0 == 1'b1 && I1 == 1'b1 && OE0 == 1'b1 && OE1 == 1'b1)
       (I2 *> ZN) = (tphlh$I2$ZN$I0_EQ_1_AN_I1_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1, tplhl$I2$ZN$I0_EQ_1_AN_I1_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1);
     if (I0 == 1'b0 && I1 == 1'b0 && OE0 == 1'b0 && OE1 == 1'b1)
       (I2 *> ZN) = (tphlh$I2$ZN$I0_EQ_0_AN_I1_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1, tplhl$I2$ZN$I0_EQ_0_AN_I1_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1);
  //   ifnone
  //     (I2 *> ZN) = (tphlh$I2$ZN,tplhl$I2$ZN);

(negedge I1 => (ZN -: ZN)) = (1.0, 1.0);

     if (I0 == 1'b1 && I2 == 1'b1 && OE0 == 1'b1 && OE1 == 1'b0)
       (I1 *> ZN) = (tphlh$I1$ZN$I0_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0, tplhl$I1$ZN$I0_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0);
     if (I0 == 1'b0 && I2 == 1'b0 && OE0 == 1'b1 && OE1 == 1'b0)
       (I1 *> ZN) = (tphlh$I1$ZN$I0_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0, tplhl$I1$ZN$I0_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0);
  //   ifnone
   //    (I1 *> ZN) = (tphlh$I1$ZN,tplhl$I1$ZN);

(negedge I0 => (ZN -: ZN)) = (1.0, 1.0);
     if (I1 == 1'b1 && I2 == 1'b1 && OE0 == 1'b0 && OE1 == 1'b0)
       (I0 *> ZN) = (tphlh$I0$ZN$I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0, tplhl$I0$ZN$I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0);
     if (I1 == 1'b0 && I2 == 1'b0 && OE0 == 1'b0 && OE1 == 1'b0)
       (I0 *> ZN) = (tphlh$I0$ZN$I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0, tplhl$I0$ZN$I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0);
 //    ifnone
  //     (I0 *> ZN) = (tphlh$I0$ZN,tplhl$I0$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_MXI3D4 (ZN, I0, I1, I2, OE0, OE1);
input  I0 ;
input  I1 ;
input  I2 ;
input  OE0 ;
input  OE1 ;
output ZN ;

   udp_mux2 (I0_out, I0, I1, OE0);
   udp_mux2 (I1_out, I0_out, I2, OE1);
   not (ZN, I1_out);

   specify
     // delay parameters
     specparam
       tplhl$I0$ZN = 1.0,
       tphlh$I0$ZN = 1.0,
       tplhl$I1$ZN = 1.0,
       tphlh$I1$ZN = 1.0,
       tplhl$I2$ZN = 1.0,
       tphlh$I2$ZN = 1.0,
       tpllh$OE0$ZN = 1.0,
       tplhl$OE0$ZN = 1.0,
       tphlh$OE0$ZN = 1.0,
       tphhl$OE0$ZN = 1.0,
       tpllh$OE1$ZN = 1.0,
       tplhl$OE1$ZN = 1.0,
       tphlh$OE1$ZN = 1.0,
       tphhl$OE1$ZN = 1.0,
       tplhl$I0$ZN$I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphlh$I0$ZN$I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tplhl$I0$ZN$I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphlh$I0$ZN$I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tplhl$I1$ZN$I0_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tphlh$I1$ZN$I0_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tplhl$I1$ZN$I0_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tphlh$I1$ZN$I0_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tplhl$I2$ZN$I0_EQ_1_AN_I1_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1 = 1.0,
       tphlh$I2$ZN$I0_EQ_1_AN_I1_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1 = 1.0,
       tplhl$I2$ZN$I0_EQ_0_AN_I1_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1 = 1.0,
       tphlh$I2$ZN$I0_EQ_0_AN_I1_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1 = 1.0,
       tpllh$OE0$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphhl$OE0$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE1_EQ_0 = 1.0,
       tpllh$OE0$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE1_EQ_0 = 1.0,
       tphhl$OE0$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE1_EQ_0 = 1.0,
       tplhl$OE0$ZN$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE1_EQ_0 = 1.0,
       tphlh$OE0$ZN$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE1_EQ_0 = 1.0,
       tplhl$OE0$ZN$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphlh$OE0$ZN$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE1_EQ_0 = 1.0,
       tpllh$OE1$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE0_EQ_1 = 1.0,
       tphhl$OE1$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE0_EQ_1 = 1.0,
       tpllh$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0 = 1.0,
       tphhl$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0 = 1.0,
       tplhl$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_1 = 1.0,
       tphlh$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_1 = 1.0,
       tplhl$OE1$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_0 = 1.0,
       tphlh$OE1$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_0 = 1.0;

     // path delays
      (posedge OE1 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge OE1 => (ZN -: ZN)) = (1.0, 1.0);
     if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && OE0 == 1'b1)
       (OE1 *> ZN) = (tpllh$OE1$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE0_EQ_1, tphhl$OE1$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE0_EQ_1);
     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && OE0 == 1'b1)
       (OE1 *> ZN) = (tphlh$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_1, tplhl$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_1);
     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && OE0 == 1'b0)
       (OE1 *> ZN) = (tpllh$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0, tphhl$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0);
     if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && OE0 == 1'b0)
       (OE1 *> ZN) = (tphlh$OE1$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_0, tplhl$OE1$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE0_EQ_0);
  //   ifnone
  //     (OE1 *> ZN) = (tpllh$OE1$ZN,tplhl$OE1$ZN);
      (posedge OE0 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge OE0 => (ZN -: ZN)) = (1.0, 1.0);
     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && OE1 == 1'b0)
       (OE0 *> ZN) = (tpllh$OE0$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE1_EQ_0, tphhl$OE0$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_OE1_EQ_0);
     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && OE1 == 1'b0)
       (OE0 *> ZN) = (tpllh$OE0$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE1_EQ_0, tphhl$OE0$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE1_EQ_0);
     if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && OE1 == 1'b0)
       (OE0 *> ZN) = (tphlh$OE0$ZN$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE1_EQ_0, tplhl$OE0$ZN$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE1_EQ_0);
     if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && OE1 == 1'b0)
       (OE0 *> ZN) = (tphlh$OE0$ZN$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE1_EQ_0, tplhl$OE0$ZN$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_OE1_EQ_0);
  //   ifnone
  //     (OE0 *> ZN) = (tpllh$OE0$ZN,tplhl$OE0$ZN);
(negedge I2 => (ZN -: ZN)) = (1.0, 1.0);
     if (I0 == 1'b1 && I1 == 1'b1 && OE0 == 1'b1 && OE1 == 1'b1)
       (I2 *> ZN) = (tphlh$I2$ZN$I0_EQ_1_AN_I1_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1, tplhl$I2$ZN$I0_EQ_1_AN_I1_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1);
     if (I0 == 1'b0 && I1 == 1'b0 && OE0 == 1'b0 && OE1 == 1'b1)
       (I2 *> ZN) = (tphlh$I2$ZN$I0_EQ_0_AN_I1_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1, tplhl$I2$ZN$I0_EQ_0_AN_I1_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1);
    // ifnone
    //   (I2 *> ZN) = (tphlh$I2$ZN,tplhl$I2$ZN);
(negedge I1 => (ZN -: ZN)) = (1.0, 1.0);
     if (I0 == 1'b1 && I2 == 1'b1 && OE0 == 1'b1 && OE1 == 1'b0)
       (I1 *> ZN) = (tphlh$I1$ZN$I0_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0, tplhl$I1$ZN$I0_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0);
     if (I0 == 1'b0 && I2 == 1'b0 && OE0 == 1'b1 && OE1 == 1'b0)
       (I1 *> ZN) = (tphlh$I1$ZN$I0_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0, tplhl$I1$ZN$I0_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0);
  //   ifnone
  //     (I1 *> ZN) = (tphlh$I1$ZN,tplhl$I1$ZN);
(negedge I0 => (ZN -: ZN)) = (1.0, 1.0);
     if (I1 == 1'b1 && I2 == 1'b1 && OE0 == 1'b0 && OE1 == 1'b0)
       (I0 *> ZN) = (tphlh$I0$ZN$I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0, tplhl$I0$ZN$I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0);
     if (I1 == 1'b0 && I2 == 1'b0 && OE0 == 1'b0 && OE1 == 1'b0)
       (I0 *> ZN) = (tphlh$I0$ZN$I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0, tplhl$I0$ZN$I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0);
 //    ifnone
 //      (I0 *> ZN) = (tphlh$I0$ZN,tplhl$I0$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_MXI4D1 (ZN, I0, I1, I2, I3, OE0, OE1);
input  I0 ;
input  I1 ;
input  I2 ;
input  I3 ;
input  OE0 ;
input  OE1 ;
output ZN ;

   udp_mux2 (I0_out, I2, I3, OE0);
   udp_mux2 (I1_out, I0, I1, OE0);
   udp_mux2 (I2_out, I1_out, I0_out, OE1);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tplhl$I0$ZN = 1.0,
       tphlh$I0$ZN = 1.0,
       tplhl$I1$ZN = 1.0,
       tphlh$I1$ZN = 1.0,
       tplhl$I2$ZN = 1.0,
       tphlh$I2$ZN = 1.0,
       tplhl$I3$ZN = 1.0,
       tphlh$I3$ZN = 1.0,
       tpllh$OE0$ZN = 1.0,
       tplhl$OE0$ZN = 1.0,
       tphlh$OE0$ZN = 1.0,
       tphhl$OE0$ZN = 1.0,
       tpllh$OE1$ZN = 1.0,
       tplhl$OE1$ZN = 1.0,
       tphlh$OE1$ZN = 1.0,
       tphhl$OE1$ZN = 1.0,
       tplhl$I0$ZN$I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphlh$I0$ZN$I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tplhl$I0$ZN$I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphlh$I0$ZN$I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tplhl$I1$ZN$I0_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tphlh$I1$ZN$I0_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tplhl$I1$ZN$I0_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tphlh$I1$ZN$I0_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tplhl$I2$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_1 = 1.0,
       tphlh$I2$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_1 = 1.0,
       tplhl$I2$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1 = 1.0,
       tphlh$I2$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1 = 1.0,
       tplhl$I3$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_1 = 1.0,
       tphlh$I3$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_1 = 1.0,
       tplhl$I3$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1 = 1.0,
       tphlh$I3$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1 = 1.0,
       tpllh$OE0$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphhl$OE0$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0 = 1.0,
       tpllh$OE0$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE1_EQ_1 = 1.0,
       tphhl$OE0$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE1_EQ_1 = 1.0,
       tplhl$OE0$ZN$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphlh$OE0$ZN$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0 = 1.0,
       tplhl$OE0$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_1_AN_OE1_EQ_1 = 1.0,
       tphlh$OE0$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_1_AN_OE1_EQ_1 = 1.0,
       tpllh$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0 = 1.0,
       tphhl$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0 = 1.0,
       tpllh$OE1$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_1 = 1.0,
       tphhl$OE1$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_1 = 1.0,
       tplhl$OE1$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_0 = 1.0,
       tphlh$OE1$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_0 = 1.0,
       tplhl$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1 = 1.0,
       tphlh$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1 = 1.0;

     // path delays
      (posedge OE1 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge OE1 => (ZN -: ZN)) = (1.0, 1.0);
     if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && OE0 == 1'b1)
       (OE1 *> ZN) = (tpllh$OE1$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_1, tphhl$OE1$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_1);
     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && OE0 == 1'b1)
       (OE1 *> ZN) = (tphlh$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1, tplhl$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1);
     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && OE0 == 1'b0)
       (OE1 *> ZN) = (tpllh$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0, tphhl$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0);
     if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && OE0 == 1'b0)
       (OE1 *> ZN) = (tphlh$OE1$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_0, tplhl$OE1$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_0);
   //  ifnone
   //    (OE1 *> ZN) = (tpllh$OE1$ZN,tplhl$OE1$ZN);
      (posedge OE0 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge OE0 => (ZN -: ZN)) = (1.0, 1.0);
     if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && OE1 == 1'b1)
       (OE0 *> ZN) = (tpllh$OE0$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE1_EQ_1, tphhl$OE0$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE1_EQ_1);
     if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && OE1 == 1'b1)
       (OE0 *> ZN) = (tphlh$OE0$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_1_AN_OE1_EQ_1, tplhl$OE0$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_1_AN_OE1_EQ_1);
     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && OE1 == 1'b0)
       (OE0 *> ZN) = (tpllh$OE0$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0, tphhl$OE0$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0);
     if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && OE1 == 1'b0)
       (OE0 *> ZN) = (tphlh$OE0$ZN$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0, tplhl$OE0$ZN$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0);
  //   ifnone
 //      (OE0 *> ZN) = (tpllh$OE0$ZN,tplhl$OE0$ZN);
(negedge I3 => (ZN -: ZN)) = (1.0, 1.0);
     if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && OE0 == 1'b1 && OE1 == 1'b1)
       (I3 *> ZN) = (tphlh$I3$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1, tplhl$I3$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1);
     if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && OE0 == 1'b1 && OE1 == 1'b1)
       (I3 *> ZN) = (tphlh$I3$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_1, tplhl$I3$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_1);
  //   ifnone
   //    (I3 *> ZN) = (tphlh$I3$ZN,tplhl$I3$ZN);
(negedge I2 => (ZN -: ZN)) = (1.0, 1.0);
     if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b1 && OE0 == 1'b0 && OE1 == 1'b1)
       (I2 *> ZN) = (tphlh$I2$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_1, tplhl$I2$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_1);
     if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b0 && OE0 == 1'b0 && OE1 == 1'b1)
       (I2 *> ZN) = (tphlh$I2$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1, tplhl$I2$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1);
  //   ifnone
    //   (I2 *> ZN) = (tphlh$I2$ZN,tplhl$I2$ZN);
(negedge I1 => (ZN -: ZN)) = (1.0, 1.0);
     if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && OE0 == 1'b1 && OE1 == 1'b0)
       (I1 *> ZN) = (tphlh$I1$ZN$I0_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0, tplhl$I1$ZN$I0_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0);
     if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && OE0 == 1'b1 && OE1 == 1'b0)
       (I1 *> ZN) = (tphlh$I1$ZN$I0_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0, tplhl$I1$ZN$I0_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0);
   //  ifnone
    //   (I1 *> ZN) = (tphlh$I1$ZN,tplhl$I1$ZN);
(negedge I0 => (ZN -: ZN)) = (1.0, 1.0);
     if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && OE0 == 1'b0 && OE1 == 1'b0)
       (I0 *> ZN) = (tphlh$I0$ZN$I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0, tplhl$I0$ZN$I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0);
     if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && OE0 == 1'b0 && OE1 == 1'b0)
       (I0 *> ZN) = (tphlh$I0$ZN$I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0, tplhl$I0$ZN$I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0);
   //  ifnone
   //    (I0 *> ZN) = (tphlh$I0$ZN,tplhl$I0$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_MXI4D2 (ZN, I0, I1, I2, I3, OE0, OE1);
input  I0 ;
input  I1 ;
input  I2 ;
input  I3 ;
input  OE0 ;
input  OE1 ;
output ZN ;

   udp_mux2 (I0_out, I2, I3, OE0);
   udp_mux2 (I1_out, I0, I1, OE0);
   udp_mux2 (I2_out, I1_out, I0_out, OE1);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tplhl$I0$ZN = 1.0,
       tphlh$I0$ZN = 1.0,
       tplhl$I1$ZN = 1.0,
       tphlh$I1$ZN = 1.0,
       tplhl$I2$ZN = 1.0,
       tphlh$I2$ZN = 1.0,
       tplhl$I3$ZN = 1.0,
       tphlh$I3$ZN = 1.0,
       tpllh$OE0$ZN = 1.0,
       tplhl$OE0$ZN = 1.0,
       tphlh$OE0$ZN = 1.0,
       tphhl$OE0$ZN = 1.0,
       tpllh$OE1$ZN = 1.0,
       tplhl$OE1$ZN = 1.0,
       tphlh$OE1$ZN = 1.0,
       tphhl$OE1$ZN = 1.0,
       tplhl$I0$ZN$I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphlh$I0$ZN$I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tplhl$I0$ZN$I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphlh$I0$ZN$I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tplhl$I1$ZN$I0_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tphlh$I1$ZN$I0_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tplhl$I1$ZN$I0_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tphlh$I1$ZN$I0_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tplhl$I2$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_1 = 1.0,
       tphlh$I2$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_1 = 1.0,
       tplhl$I2$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1 = 1.0,
       tphlh$I2$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1 = 1.0,
       tplhl$I3$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_1 = 1.0,
       tphlh$I3$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_1 = 1.0,
       tplhl$I3$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1 = 1.0,
       tphlh$I3$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1 = 1.0,
       tpllh$OE0$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphhl$OE0$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0 = 1.0,
       tpllh$OE0$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE1_EQ_1 = 1.0,
       tphhl$OE0$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE1_EQ_1 = 1.0,
       tplhl$OE0$ZN$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphlh$OE0$ZN$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0 = 1.0,
       tplhl$OE0$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_1_AN_OE1_EQ_1 = 1.0,
       tphlh$OE0$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_1_AN_OE1_EQ_1 = 1.0,
       tpllh$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0 = 1.0,
       tphhl$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0 = 1.0,
       tpllh$OE1$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_1 = 1.0,
       tphhl$OE1$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_1 = 1.0,
       tplhl$OE1$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_0 = 1.0,
       tphlh$OE1$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_0 = 1.0,
       tplhl$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1 = 1.0,
       tphlh$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1 = 1.0;

     // path delays
      (posedge OE1 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge OE1 => (ZN -: ZN)) = (1.0, 1.0);

     if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && OE0 == 1'b1)
       (OE1 *> ZN) = (tpllh$OE1$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_1, tphhl$OE1$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_1);
     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && OE0 == 1'b1)
       (OE1 *> ZN) = (tphlh$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1, tplhl$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1);
     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && OE0 == 1'b0)
       (OE1 *> ZN) = (tpllh$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0, tphhl$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0);
     if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && OE0 == 1'b0)
       (OE1 *> ZN) = (tphlh$OE1$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_0, tplhl$OE1$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_0);
   //  ifnone
    //   (OE1 *> ZN) = (tpllh$OE1$ZN,tplhl$OE1$ZN);

      (posedge OE0 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge OE0 => (ZN -: ZN)) = (1.0, 1.0);

     if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && OE1 == 1'b1)
       (OE0 *> ZN) = (tpllh$OE0$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE1_EQ_1, tphhl$OE0$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE1_EQ_1);
     if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && OE1 == 1'b1)
       (OE0 *> ZN) = (tphlh$OE0$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_1_AN_OE1_EQ_1, tplhl$OE0$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_1_AN_OE1_EQ_1);
     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && OE1 == 1'b0)
       (OE0 *> ZN) = (tpllh$OE0$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0, tphhl$OE0$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0);
     if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && OE1 == 1'b0)
       (OE0 *> ZN) = (tphlh$OE0$ZN$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0, tplhl$OE0$ZN$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0);
   //  ifnone
   //    (OE0 *> ZN) = (tpllh$OE0$ZN,tplhl$OE0$ZN);
(negedge I3 => (ZN -: ZN)) = (1.0, 1.0);
     if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && OE0 == 1'b1 && OE1 == 1'b1)
       (I3 *> ZN) = (tphlh$I3$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1, tplhl$I3$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1);
     if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && OE0 == 1'b1 && OE1 == 1'b1)
       (I3 *> ZN) = (tphlh$I3$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_1, tplhl$I3$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_1);
   //  ifnone
   //    (I3 *> ZN) = (tphlh$I3$ZN,tplhl$I3$ZN);
(negedge I2 => (ZN -: ZN)) = (1.0, 1.0);
     if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b1 && OE0 == 1'b0 && OE1 == 1'b1)
       (I2 *> ZN) = (tphlh$I2$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_1, tplhl$I2$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_1);
     if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b0 && OE0 == 1'b0 && OE1 == 1'b1)
       (I2 *> ZN) = (tphlh$I2$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1, tplhl$I2$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1);
   //  ifnone
  //     (I2 *> ZN) = (tphlh$I2$ZN,tplhl$I2$ZN);
(negedge I1 => (ZN -: ZN)) = (1.0, 1.0);
     if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && OE0 == 1'b1 && OE1 == 1'b0)
       (I1 *> ZN) = (tphlh$I1$ZN$I0_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0, tplhl$I1$ZN$I0_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0);
     if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && OE0 == 1'b1 && OE1 == 1'b0)
       (I1 *> ZN) = (tphlh$I1$ZN$I0_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0, tplhl$I1$ZN$I0_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0);
 //    ifnone
  //     (I1 *> ZN) = (tphlh$I1$ZN,tplhl$I1$ZN);
(negedge I0 => (ZN -: ZN)) = (1.0, 1.0);
     if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && OE0 == 1'b0 && OE1 == 1'b0)
       (I0 *> ZN) = (tphlh$I0$ZN$I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0, tplhl$I0$ZN$I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0);
     if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && OE0 == 1'b0 && OE1 == 1'b0)
       (I0 *> ZN) = (tphlh$I0$ZN$I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0, tplhl$I0$ZN$I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0);
 //    ifnone
//       (I0 *> ZN) = (tphlh$I0$ZN,tplhl$I0$ZN);
//



   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_MXI4D4 (ZN, I0, I1, I2, I3, OE0, OE1);
input  I0 ;
input  I1 ;
input  I2 ;
input  I3 ;
input  OE0 ;
input  OE1 ;
output ZN ;

   udp_mux2 (I0_out, I2, I3, OE0);
   udp_mux2 (I1_out, I0, I1, OE0);
   udp_mux2 (I2_out, I1_out, I0_out, OE1);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tplhl$I0$ZN = 1.0,
       tphlh$I0$ZN = 1.0,
       tplhl$I1$ZN = 1.0,
       tphlh$I1$ZN = 1.0,
       tplhl$I2$ZN = 1.0,
       tphlh$I2$ZN = 1.0,
       tplhl$I3$ZN = 1.0,
       tphlh$I3$ZN = 1.0,
       tpllh$OE0$ZN = 1.0,
       tplhl$OE0$ZN = 1.0,
       tphlh$OE0$ZN = 1.0,
       tphhl$OE0$ZN = 1.0,
       tpllh$OE1$ZN = 1.0,
       tplhl$OE1$ZN = 1.0,
       tphlh$OE1$ZN = 1.0,
       tphhl$OE1$ZN = 1.0,
       tplhl$I0$ZN$I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphlh$I0$ZN$I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tplhl$I0$ZN$I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphlh$I0$ZN$I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0 = 1.0,
       tplhl$I1$ZN$I0_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tphlh$I1$ZN$I0_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tplhl$I1$ZN$I0_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tphlh$I1$ZN$I0_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0 = 1.0,
       tplhl$I2$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_1 = 1.0,
       tphlh$I2$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_1 = 1.0,
       tplhl$I2$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1 = 1.0,
       tphlh$I2$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1 = 1.0,
       tplhl$I3$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_1 = 1.0,
       tphlh$I3$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_1 = 1.0,
       tplhl$I3$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1 = 1.0,
       tphlh$I3$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1 = 1.0,
       tpllh$OE0$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphhl$OE0$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0 = 1.0,
       tpllh$OE0$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE1_EQ_1 = 1.0,
       tphhl$OE0$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE1_EQ_1 = 1.0,
       tplhl$OE0$ZN$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0 = 1.0,
       tphlh$OE0$ZN$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0 = 1.0,
       tplhl$OE0$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_1_AN_OE1_EQ_1 = 1.0,
       tphlh$OE0$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_1_AN_OE1_EQ_1 = 1.0,
       tpllh$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0 = 1.0,
       tphhl$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0 = 1.0,
       tpllh$OE1$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_1 = 1.0,
       tphhl$OE1$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_1 = 1.0,
       tplhl$OE1$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_0 = 1.0,
       tphlh$OE1$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_0 = 1.0,
       tplhl$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1 = 1.0,
       tphlh$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1 = 1.0;

     // path delays
      (posedge OE1 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge OE1 => (ZN -: ZN)) = (1.0, 1.0);

     if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && OE0 == 1'b1)
       (OE1 *> ZN) = (tpllh$OE1$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_1, tphhl$OE1$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_1);
     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && OE0 == 1'b1)
       (OE1 *> ZN) = (tphlh$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1, tplhl$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1);
     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && OE0 == 1'b0)
       (OE1 *> ZN) = (tpllh$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0, tphhl$OE1$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0);
     if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && OE0 == 1'b0)
       (OE1 *> ZN) = (tphlh$OE1$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_0, tplhl$OE1$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE0_EQ_0);
 //    ifnone
   //    (OE1 *> ZN) = (tpllh$OE1$ZN,tplhl$OE1$ZN);
      (posedge OE0 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge OE0 => (ZN -: ZN)) = (1.0, 1.0);
     if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && OE1 == 1'b1)
       (OE0 *> ZN) = (tpllh$OE0$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE1_EQ_1, tphhl$OE0$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_0_AN_OE1_EQ_1);
     if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && OE1 == 1'b1)
       (OE0 *> ZN) = (tphlh$OE0$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_1_AN_OE1_EQ_1, tplhl$OE0$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_1_AN_OE1_EQ_1);
     if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && OE1 == 1'b0)
       (OE0 *> ZN) = (tpllh$OE0$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0, tphhl$OE0$ZN$I0_EQ_1_AN_I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0);
     if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && OE1 == 1'b0)
       (OE0 *> ZN) = (tphlh$OE0$ZN$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0, tplhl$OE0$ZN$I0_EQ_0_AN_I1_EQ_1_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE1_EQ_0);
   //  ifnone
     //  (OE0 *> ZN) = (tpllh$OE0$ZN,tplhl$OE0$ZN);
      (negedge I3 => (ZN -: ZN)) = (1.0, 1.0);
     if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && OE0 == 1'b1 && OE1 == 1'b1)
       (I3 *> ZN) = (tphlh$I3$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1, tplhl$I3$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I2_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_1);
     if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && OE0 == 1'b1 && OE1 == 1'b1)
       (I3 *> ZN) = (tphlh$I3$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_1, tplhl$I3$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I2_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_1);
   //  ifnone
     //  (I3 *> ZN) = (tphlh$I3$ZN,tplhl$I3$ZN);

(negedge I2 => (ZN -: ZN)) = (1.0, 1.0);
     if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b1 && OE0 == 1'b0 && OE1 == 1'b1)
       (I2 *> ZN) = (tphlh$I2$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_1, tplhl$I2$ZN$I0_EQ_1_AN_I1_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_1);
     if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b0 && OE0 == 1'b0 && OE1 == 1'b1)
       (I2 *> ZN) = (tphlh$I2$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1, tplhl$I2$ZN$I0_EQ_0_AN_I1_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_1);
  ///   ifnone
    //   (I2 *> ZN) = (tphlh$I2$ZN,tplhl$I2$ZN);

(negedge I1 => (ZN -: ZN)) = (1.0, 1.0);
     if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && OE0 == 1'b1 && OE1 == 1'b0)
       (I1 *> ZN) = (tphlh$I1$ZN$I0_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0, tplhl$I1$ZN$I0_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_1_AN_OE1_EQ_0);
     if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && OE0 == 1'b1 && OE1 == 1'b0)
       (I1 *> ZN) = (tphlh$I1$ZN$I0_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0, tplhl$I1$ZN$I0_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_1_AN_OE1_EQ_0);
  //   ifnone
  //     (I1 *> ZN) = (tphlh$I1$ZN,tplhl$I1$ZN);

(negedge I0 => (ZN -: ZN)) = (1.0, 1.0);
     if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && OE0 == 1'b0 && OE1 == 1'b0)
       (I0 *> ZN) = (tphlh$I0$ZN$I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0, tplhl$I0$ZN$I1_EQ_1_AN_I2_EQ_1_AN_I3_EQ_1_AN_OE0_EQ_0_AN_OE1_EQ_0);
     if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && OE0 == 1'b0 && OE1 == 1'b0)
       (I0 *> ZN) = (tphlh$I0$ZN$I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0, tplhl$I0$ZN$I1_EQ_0_AN_I2_EQ_0_AN_I3_EQ_0_AN_OE0_EQ_0_AN_OE1_EQ_0);
  //   ifnone
  //     (I0 *> ZN) = (tphlh$I0$ZN,tplhl$I0$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_ND02BD1 (ZN, A1N, A2);
input  A1N ;
input  A2 ;
output ZN ;

   not (I0_out, A1N);
   and (I1_out, I0_out, A2);
   not (ZN, I1_out);

   specify
     // delay parameters
     specparam
       tpllh$A1N$ZN = 1.0,
       tphhl$A1N$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0;

     // path delays
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1N *> ZN) = (tpllh$A1N$ZN, tphhl$A1N$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_ND02BD2 (ZN, A1N, A2);
input  A1N ;
input  A2 ;
output ZN ;

   not (I0_out, A1N);
   and (I1_out, I0_out, A2);
   not (ZN, I1_out);

   specify
     // delay parameters
     specparam
       tpllh$A1N$ZN = 1.0,
       tphhl$A1N$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0;

     // path delays
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1N *> ZN) = (tpllh$A1N$ZN, tphhl$A1N$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_ND02BD4 (ZN, A1N, A2);
input  A1N ;
input  A2 ;
output ZN ;

   not (I0_out, A1N);
   and (I1_out, I0_out, A2);
   not (ZN, I1_out);

   specify
     // delay parameters
     specparam
       tpllh$A1N$ZN = 1.0,
       tphhl$A1N$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0;

     // path delays
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1N *> ZN) = (tpllh$A1N$ZN, tphhl$A1N$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_ND02D1 (ZN, A1, A2);
input  A1 ;
input  A2 ;
output ZN ;

   and (I0_out, A1, A2);
   not (ZN, I0_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0;

     // path delays
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_ND02D2 (ZN, A1, A2);
input  A1 ;
input  A2 ;
output ZN ;

   and (I0_out, A1, A2);
   not (ZN, I0_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0;

     // path delays
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_ND02D4 (ZN, A1, A2);
input  A1 ;
input  A2 ;
output ZN ;

   and (I0_out, A1, A2);
   not (ZN, I0_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0;

     // path delays
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_ND03BD1 (ZN, A1N, A2, A3);
input  A1N ;
input  A2 ;
input  A3 ;
output ZN ;

   not (I0_out, A1N);
   and (I2_out, I0_out, A2, A3);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tpllh$A1N$ZN = 1.0,
       tphhl$A1N$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0;

     // path delays
     (A3 *> ZN) = (tphlh$A3$ZN, tplhl$A3$ZN);
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1N *> ZN) = (tpllh$A1N$ZN, tphhl$A1N$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_ND03BD2 (ZN, A1N, A2, A3);
input  A1N ;
input  A2 ;
input  A3 ;
output ZN ;

   not (I0_out, A1N);
   and (I2_out, I0_out, A2, A3);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tpllh$A1N$ZN = 1.0,
       tphhl$A1N$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0;

     // path delays
     (A3 *> ZN) = (tphlh$A3$ZN, tplhl$A3$ZN);
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1N *> ZN) = (tpllh$A1N$ZN, tphhl$A1N$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_ND03BD4 (ZN, A1N, A2, A3);
input  A1N ;
input  A2 ;
input  A3 ;
output ZN ;

   not (I0_out, A1N);
   and (I2_out, I0_out, A2, A3);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tpllh$A1N$ZN = 1.0,
       tphhl$A1N$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0;

     // path delays
     (A3 *> ZN) = (tphlh$A3$ZN, tplhl$A3$ZN);
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1N *> ZN) = (tpllh$A1N$ZN, tphhl$A1N$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_ND03D1 (ZN, A1, A2, A3);
input  A1 ;
input  A2 ;
input  A3 ;
output ZN ;

   and (I1_out, A1, A2, A3);
   not (ZN, I1_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0;

     // path delays
     (A3 *> ZN) = (tphlh$A3$ZN, tplhl$A3$ZN);
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_ND03D2 (ZN, A1, A2, A3);
input  A1 ;
input  A2 ;
input  A3 ;
output ZN ;

   and (I1_out, A1, A2, A3);
   not (ZN, I1_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0;

     // path delays
     (A3 *> ZN) = (tphlh$A3$ZN, tplhl$A3$ZN);
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_ND03D4 (ZN, A1, A2, A3);
input  A1 ;
input  A2 ;
input  A3 ;
output ZN ;

   and (I1_out, A1, A2, A3);
   not (ZN, I1_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0;

     // path delays
     (A3 *> ZN) = (tphlh$A3$ZN, tplhl$A3$ZN);
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_ND04BBD1 (ZN, A1N, A2N, A3, A4);
input  A1N ;
input  A2N ;
input  A3 ;
input  A4 ;
output ZN ;

   not (I0_out, A1N);
   not (I1_out, A2N);
   and (I4_out, I0_out, I1_out, A3, A4);
   not (ZN, I4_out);

   specify
     // delay parameters
     specparam
       tpllh$A1N$ZN = 1.0,
       tphhl$A1N$ZN = 1.0,
       tpllh$A2N$ZN = 1.0,
       tphhl$A2N$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0,
       tplhl$A4$ZN = 1.0,
       tphlh$A4$ZN = 1.0;

     // path delays
     (A4 *> ZN) = (tphlh$A4$ZN, tplhl$A4$ZN);
     (A3 *> ZN) = (tphlh$A3$ZN, tplhl$A3$ZN);
     (A2N *> ZN) = (tpllh$A2N$ZN, tphhl$A2N$ZN);
     (A1N *> ZN) = (tpllh$A1N$ZN, tphhl$A1N$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_ND04BBD2 (ZN, A1N, A2N, A3, A4);
input  A1N ;
input  A2N ;
input  A3 ;
input  A4 ;
output ZN ;

   not (I0_out, A1N);
   not (I1_out, A2N);
   and (I4_out, I0_out, I1_out, A3, A4);
   not (ZN, I4_out);

   specify
     // delay parameters
     specparam
       tpllh$A1N$ZN = 1.0,
       tphhl$A1N$ZN = 1.0,
       tpllh$A2N$ZN = 1.0,
       tphhl$A2N$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0,
       tplhl$A4$ZN = 1.0,
       tphlh$A4$ZN = 1.0;

     // path delays
     (A4 *> ZN) = (tphlh$A4$ZN, tplhl$A4$ZN);
     (A3 *> ZN) = (tphlh$A3$ZN, tplhl$A3$ZN);
     (A2N *> ZN) = (tpllh$A2N$ZN, tphhl$A2N$ZN);
     (A1N *> ZN) = (tpllh$A1N$ZN, tphhl$A1N$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_ND04BBD4 (ZN, A1N, A2N, A3, A4);
input  A1N ;
input  A2N ;
input  A3 ;
input  A4 ;
output ZN ;

   not (I0_out, A2N);
   not (I1_out, A1N);
   and (I4_out, I0_out, I1_out, A3, A4);
   not (ZN, I4_out);

   specify
     // delay parameters
     specparam
       tpllh$A1N$ZN = 1.0,
       tphhl$A1N$ZN = 1.0,
       tpllh$A2N$ZN = 1.0,
       tphhl$A2N$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0,
       tplhl$A4$ZN = 1.0,
       tphlh$A4$ZN = 1.0;

     // path delays
     (A4 *> ZN) = (tphlh$A4$ZN, tplhl$A4$ZN);
     (A3 *> ZN) = (tphlh$A3$ZN, tplhl$A3$ZN);
     (A2N *> ZN) = (tpllh$A2N$ZN, tphhl$A2N$ZN);
     (A1N *> ZN) = (tpllh$A1N$ZN, tphhl$A1N$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_ND04BD1 (ZN, A1N, A2, A3, A4);
input  A1N ;
input  A2 ;
input  A3 ;
input  A4 ;
output ZN ;

   not (I0_out, A1N);
   and (I3_out, I0_out, A2, A3, A4);
   not (ZN, I3_out);

   specify
     // delay parameters
     specparam
       tpllh$A1N$ZN = 1.0,
       tphhl$A1N$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0,
       tplhl$A4$ZN = 1.0,
       tphlh$A4$ZN = 1.0;

     // path delays
     (A4 *> ZN) = (tphlh$A4$ZN, tplhl$A4$ZN);
     (A3 *> ZN) = (tphlh$A3$ZN, tplhl$A3$ZN);
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1N *> ZN) = (tpllh$A1N$ZN, tphhl$A1N$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_ND04BD2 (ZN, A1N, A2, A3, A4);
input  A1N ;
input  A2 ;
input  A3 ;
input  A4 ;
output ZN ;

   not (I0_out, A1N);
   and (I3_out, I0_out, A2, A3, A4);
   not (ZN, I3_out);

   specify
     // delay parameters
     specparam
       tpllh$A1N$ZN = 1.0,
       tphhl$A1N$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0,
       tplhl$A4$ZN = 1.0,
       tphlh$A4$ZN = 1.0;

     // path delays
     (A4 *> ZN) = (tphlh$A4$ZN, tplhl$A4$ZN);
     (A3 *> ZN) = (tphlh$A3$ZN, tplhl$A3$ZN);
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1N *> ZN) = (tpllh$A1N$ZN, tphhl$A1N$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_ND04BD4 (ZN, A1N, A2, A3, A4);
input  A1N ;
input  A2 ;
input  A3 ;
input  A4 ;
output ZN ;

   not (I0_out, A1N);
   and (I3_out, I0_out, A2, A3, A4);
   not (ZN, I3_out);

   specify
     // delay parameters
     specparam
       tpllh$A1N$ZN = 1.0,
       tphhl$A1N$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0,
       tplhl$A4$ZN = 1.0,
       tphlh$A4$ZN = 1.0;

     // path delays
     (A4 *> ZN) = (tphlh$A4$ZN, tplhl$A4$ZN);
     (A3 *> ZN) = (tphlh$A3$ZN, tplhl$A3$ZN);
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1N *> ZN) = (tpllh$A1N$ZN, tphhl$A1N$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_ND04D1 (ZN, A1, A2, A3, A4);
input  A1 ;
input  A2 ;
input  A3 ;
input  A4 ;
output ZN ;

   and (I2_out, A1, A2, A3, A4);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0,
       tplhl$A4$ZN = 1.0,
       tphlh$A4$ZN = 1.0;

     // path delays
     (A4 *> ZN) = (tphlh$A4$ZN, tplhl$A4$ZN);
     (A3 *> ZN) = (tphlh$A3$ZN, tplhl$A3$ZN);
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_ND04D2 (ZN, A1, A2, A3, A4);
input  A1 ;
input  A2 ;
input  A3 ;
input  A4 ;
output ZN ;

   and (I2_out, A1, A2, A3, A4);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0,
       tplhl$A4$ZN = 1.0,
       tphlh$A4$ZN = 1.0;

     // path delays
     (A4 *> ZN) = (tphlh$A4$ZN, tplhl$A4$ZN);
     (A3 *> ZN) = (tphlh$A3$ZN, tplhl$A3$ZN);
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_ND04D4 (ZN, A1, A2, A3, A4);
input  A1 ;
input  A2 ;
input  A3 ;
input  A4 ;
output ZN ;

   and (I2_out, A1, A2, A3, A4);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0,
       tplhl$A4$ZN = 1.0,
       tphlh$A4$ZN = 1.0;

     // path delays
     (A4 *> ZN) = (tphlh$A4$ZN, tplhl$A4$ZN);
     (A3 *> ZN) = (tphlh$A3$ZN, tplhl$A3$ZN);
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_NR02BD1 (ZN, A1N, A2);
input  A1N ;
input  A2 ;
output ZN ;

   not (I0_out, A1N);
   or  (I1_out, I0_out, A2);
   not (ZN, I1_out);

   specify
     // delay parameters
     specparam
       tpllh$A1N$ZN = 1.0,
       tphhl$A1N$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0;

     // path delays
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1N *> ZN) = (tpllh$A1N$ZN, tphhl$A1N$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_NR02BD2 (ZN, A1N, A2);
input  A1N ;
input  A2 ;
output ZN ;

   not (I0_out, A1N);
   or  (I1_out, I0_out, A2);
   not (ZN, I1_out);

   specify
     // delay parameters
     specparam
       tpllh$A1N$ZN = 1.0,
       tphhl$A1N$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0;

     // path delays
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1N *> ZN) = (tpllh$A1N$ZN, tphhl$A1N$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_NR02BD4 (ZN, A1N, A2);
input  A1N ;
input  A2 ;
output ZN ;

   not (I0_out, A1N);
   or  (I1_out, I0_out, A2);
   not (ZN, I1_out);

   specify
     // delay parameters
     specparam
       tpllh$A1N$ZN = 1.0,
       tphhl$A1N$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0;

     // path delays
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1N *> ZN) = (tpllh$A1N$ZN, tphhl$A1N$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_NR02D1 (ZN, A1, A2);
input  A1 ;
input  A2 ;
output ZN ;

   or  (I0_out, A1, A2);
   not (ZN, I0_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0;

     // path delays
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_NR02D2 (ZN, A1, A2);
input  A1 ;
input  A2 ;
output ZN ;

   or  (I0_out, A1, A2);
   not (ZN, I0_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0;

     // path delays
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_NR02D4 (ZN, A1, A2);
input  A1 ;
input  A2 ;
output ZN ;

   or  (I0_out, A1, A2);
   not (ZN, I0_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0;

     // path delays
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_NR03BD1 (ZN, A1N, A2, A3);
input  A1N ;
input  A2 ;
input  A3 ;
output ZN ;

   not (I0_out, A1N);
   or  (I2_out, I0_out, A2, A3);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tpllh$A1N$ZN = 1.0,
       tphhl$A1N$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0;

     // path delays
     (A3 *> ZN) = (tphlh$A3$ZN, tplhl$A3$ZN);
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1N *> ZN) = (tpllh$A1N$ZN, tphhl$A1N$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_NR03BD2 (ZN, A1N, A2, A3);
input  A1N ;
input  A2 ;
input  A3 ;
output ZN ;

   not (I0_out, A1N);
   or  (I2_out, I0_out, A2, A3);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tpllh$A1N$ZN = 1.0,
       tphhl$A1N$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0;

     // path delays
     (A3 *> ZN) = (tphlh$A3$ZN, tplhl$A3$ZN);
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1N *> ZN) = (tpllh$A1N$ZN, tphhl$A1N$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_NR03BD4 (ZN, A1N, A2, A3);
input  A1N ;
input  A2 ;
input  A3 ;
output ZN ;

   not (I0_out, A1N);
   or  (I2_out, I0_out, A2, A3);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tpllh$A1N$ZN = 1.0,
       tphhl$A1N$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0;

     // path delays
     (A3 *> ZN) = (tphlh$A3$ZN, tplhl$A3$ZN);
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1N *> ZN) = (tpllh$A1N$ZN, tphhl$A1N$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_NR03D1 (ZN, A1, A2, A3);
input  A1 ;
input  A2 ;
input  A3 ;
output ZN ;

   or  (I1_out, A1, A2, A3);
   not (ZN, I1_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0;

     // path delays
     (A3 *> ZN) = (tphlh$A3$ZN, tplhl$A3$ZN);
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_NR03D2 (ZN, A1, A2, A3);
input  A1 ;
input  A2 ;
input  A3 ;
output ZN ;

   or  (I1_out, A1, A2, A3);
   not (ZN, I1_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0;

     // path delays
     (A3 *> ZN) = (tphlh$A3$ZN, tplhl$A3$ZN);
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_NR03D4 (ZN, A1, A2, A3);
input  A1 ;
input  A2 ;
input  A3 ;
output ZN ;

   or  (I1_out, A1, A2, A3);
   not (ZN, I1_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0;

     // path delays
     (A3 *> ZN) = (tphlh$A3$ZN, tplhl$A3$ZN);
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_NR04BBD1 (ZN, A1N, A2N, A3, A4);
input  A1N ;
input  A2N ;
input  A3 ;
input  A4 ;
output ZN ;

   not (I0_out, A2N);
   not (I1_out, A1N);
   or  (I4_out, I0_out, I1_out, A3, A4);
   not (ZN, I4_out);

   specify
     // delay parameters
     specparam
       tpllh$A1N$ZN = 1.0,
       tphhl$A1N$ZN = 1.0,
       tpllh$A2N$ZN = 1.0,
       tphhl$A2N$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0,
       tplhl$A4$ZN = 1.0,
       tphlh$A4$ZN = 1.0;

     // path delays
     (A4 *> ZN) = (tphlh$A4$ZN, tplhl$A4$ZN);
     (A3 *> ZN) = (tphlh$A3$ZN, tplhl$A3$ZN);
     (A2N *> ZN) = (tpllh$A2N$ZN, tphhl$A2N$ZN);
     (A1N *> ZN) = (tpllh$A1N$ZN, tphhl$A1N$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_NR04BBD2 (ZN, A1N, A2N, A3, A4);
input  A1N ;
input  A2N ;
input  A3 ;
input  A4 ;
output ZN ;

   not (I0_out, A1N);
   not (I1_out, A2N);
   or  (I4_out, I0_out, I1_out, A3, A4);
   not (ZN, I4_out);

   specify
     // delay parameters
     specparam
       tpllh$A1N$ZN = 1.0,
       tphhl$A1N$ZN = 1.0,
       tpllh$A2N$ZN = 1.0,
       tphhl$A2N$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0,
       tplhl$A4$ZN = 1.0,
       tphlh$A4$ZN = 1.0;

     // path delays
     (A4 *> ZN) = (tphlh$A4$ZN, tplhl$A4$ZN);
     (A3 *> ZN) = (tphlh$A3$ZN, tplhl$A3$ZN);
     (A2N *> ZN) = (tpllh$A2N$ZN, tphhl$A2N$ZN);
     (A1N *> ZN) = (tpllh$A1N$ZN, tphhl$A1N$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_NR04BBD4 (ZN, A1N, A2N, A3, A4);
input  A1N ;
input  A2N ;
input  A3 ;
input  A4 ;
output ZN ;

   not (I0_out, A1N);
   not (I1_out, A2N);
   or  (I4_out, I0_out, I1_out, A3, A4);
   not (ZN, I4_out);

   specify
     // delay parameters
     specparam
       tpllh$A1N$ZN = 1.0,
       tphhl$A1N$ZN = 1.0,
       tpllh$A2N$ZN = 1.0,
       tphhl$A2N$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0,
       tplhl$A4$ZN = 1.0,
       tphlh$A4$ZN = 1.0;

     // path delays
     (A4 *> ZN) = (tphlh$A4$ZN, tplhl$A4$ZN);
     (A3 *> ZN) = (tphlh$A3$ZN, tplhl$A3$ZN);
     (A2N *> ZN) = (tpllh$A2N$ZN, tphhl$A2N$ZN);
     (A1N *> ZN) = (tpllh$A1N$ZN, tphhl$A1N$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_NR04BD1 (ZN, A1N, A2, A3, A4);
input  A1N ;
input  A2 ;
input  A3 ;
input  A4 ;
output ZN ;

   not (I0_out, A1N);
   or  (I3_out, I0_out, A2, A3, A4);
   not (ZN, I3_out);

   specify
     // delay parameters
     specparam
       tpllh$A1N$ZN = 1.0,
       tphhl$A1N$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0,
       tplhl$A4$ZN = 1.0,
       tphlh$A4$ZN = 1.0;

     // path delays
     (A4 *> ZN) = (tphlh$A4$ZN, tplhl$A4$ZN);
     (A3 *> ZN) = (tphlh$A3$ZN, tplhl$A3$ZN);
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1N *> ZN) = (tpllh$A1N$ZN, tphhl$A1N$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_NR04BD2 (ZN, A1N, A2, A3, A4);
input  A1N ;
input  A2 ;
input  A3 ;
input  A4 ;
output ZN ;

   not (I0_out, A1N);
   or  (I3_out, I0_out, A2, A3, A4);
   not (ZN, I3_out);

   specify
     // delay parameters
     specparam
       tpllh$A1N$ZN = 1.0,
       tphhl$A1N$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0,
       tplhl$A4$ZN = 1.0,
       tphlh$A4$ZN = 1.0;

     // path delays
     (A4 *> ZN) = (tphlh$A4$ZN, tplhl$A4$ZN);
     (A3 *> ZN) = (tphlh$A3$ZN, tplhl$A3$ZN);
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1N *> ZN) = (tpllh$A1N$ZN, tphhl$A1N$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_NR04BD4 (ZN, A1N, A2, A3, A4);
input  A1N ;
input  A2 ;
input  A3 ;
input  A4 ;
output ZN ;

   not (I0_out, A1N);
   or  (I3_out, I0_out, A2, A3, A4);
   not (ZN, I3_out);

   specify
     // delay parameters
     specparam
       tpllh$A1N$ZN = 1.0,
       tphhl$A1N$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0,
       tplhl$A4$ZN = 1.0,
       tphlh$A4$ZN = 1.0;

     // path delays
     (A4 *> ZN) = (tphlh$A4$ZN, tplhl$A4$ZN);
     (A3 *> ZN) = (tphlh$A3$ZN, tplhl$A3$ZN);
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1N *> ZN) = (tpllh$A1N$ZN, tphhl$A1N$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_NR04D1 (ZN, A1, A2, A3, A4);
input  A1 ;
input  A2 ;
input  A3 ;
input  A4 ;
output ZN ;

   or  (I2_out, A1, A2, A3, A4);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0,
       tplhl$A4$ZN = 1.0,
       tphlh$A4$ZN = 1.0;

     // path delays
     (A4 *> ZN) = (tphlh$A4$ZN, tplhl$A4$ZN);
     (A3 *> ZN) = (tphlh$A3$ZN, tplhl$A3$ZN);
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_NR04D2 (ZN, A1, A2, A3, A4);
input  A1 ;
input  A2 ;
input  A3 ;
input  A4 ;
output ZN ;

   or  (I2_out, A1, A2, A3, A4);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0,
       tplhl$A4$ZN = 1.0,
       tphlh$A4$ZN = 1.0;

     // path delays
     (A4 *> ZN) = (tphlh$A4$ZN, tplhl$A4$ZN);
     (A3 *> ZN) = (tphlh$A3$ZN, tplhl$A3$ZN);
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_NR04D4 (ZN, A1, A2, A3, A4);
input  A1 ;
input  A2 ;
input  A3 ;
input  A4 ;
output ZN ;

   or  (I2_out, A1, A2, A3, A4);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0,
       tplhl$A4$ZN = 1.0,
       tphlh$A4$ZN = 1.0;

     // path delays
     (A4 *> ZN) = (tphlh$A4$ZN, tplhl$A4$ZN);
     (A3 *> ZN) = (tphlh$A3$ZN, tplhl$A3$ZN);
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_NT01D1 (Z, I, OE);
input  I ;
input  OE ;
output Z ;

   bufif1 (Z, I, OE);

   specify
     // delay parameters
     specparam
       tpllh$I$Z = 1.0,
       tphhl$I$Z = 1.0,
       tpzh$OE$Z = 1.0,
       tpzl$OE$Z = 1.0,
       tplz$OE$Z = 1.0,
       tphz$OE$Z = 1.0;

     // path delays
     (OE *> Z) = (0, 0, tplz$OE$Z, tpzh$OE$Z, tphz$OE$Z, tpzl$OE$Z);
     (I *> Z) = (tpllh$I$Z, tphhl$I$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_NT01D2 (Z, I, OE);
input  I ;
input  OE ;
output Z ;

   bufif1 (Z, I, OE);

   specify
     // delay parameters
     specparam
       tpllh$I$Z = 1.0,
       tphhl$I$Z = 1.0,
       tpzh$OE$Z = 1.0,
       tpzl$OE$Z = 1.0,
       tplz$OE$Z = 1.0,
       tphz$OE$Z = 1.0;

     // path delays
     (OE *> Z) = (0, 0, tplz$OE$Z, tpzh$OE$Z, tphz$OE$Z, tpzl$OE$Z);
     (I *> Z) = (tpllh$I$Z, tphhl$I$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_NT01D4 (Z, I, OE);
input  I ;
input  OE ;
output Z ;

   bufif1 (Z, I, OE);

   specify
     // delay parameters
     specparam
       tpllh$I$Z = 1.0,
       tphhl$I$Z = 1.0,
       tpzh$OE$Z = 1.0,
       tpzl$OE$Z = 1.0,
       tplz$OE$Z = 1.0,
       tphz$OE$Z = 1.0;

     // path delays
     (OE *> Z) = (0, 0, tplz$OE$Z, tpzh$OE$Z, tphz$OE$Z, tpzl$OE$Z);
     (I *> Z) = (tpllh$I$Z, tphhl$I$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_NT01D6 (Z, I, OE);
input  I ;
input  OE ;
output Z ;

   bufif1 (Z, I, OE);

   specify
     // delay parameters
     specparam
       tpllh$I$Z = 1.0,
       tphhl$I$Z = 1.0,
       tpzh$OE$Z = 1.0,
       tpzl$OE$Z = 1.0,
       tplz$OE$Z = 1.0,
       tphz$OE$Z = 1.0;

     // path delays
     (OE *> Z) = (0, 0, tplz$OE$Z, tpzh$OE$Z, tphz$OE$Z, tpzl$OE$Z);
     (I *> Z) = (tpllh$I$Z, tphhl$I$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_NT02D1 (Z, I, OE);
input  I ;
input  OE ;
output Z ;

   bufif0 (Z, I, OE);

   specify
     // delay parameters
     specparam
       tpllh$I$Z = 1.0,
       tphhl$I$Z = 1.0,
       tplz$OE$Z = 1.0,
       tphz$OE$Z = 1.0,
       tpzh$OE$Z = 1.0,
       tpzl$OE$Z = 1.0;

     // path delays
     (OE *> Z) = (0, 0, tplz$OE$Z, tpzh$OE$Z, tphz$OE$Z, tpzl$OE$Z);
     (I *> Z) = (tpllh$I$Z, tphhl$I$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_NT02D2 (Z, I, OE);
input  I ;
input  OE ;
output Z ;

   bufif0 (Z, I, OE);

   specify
     // delay parameters
     specparam
       tpllh$I$Z = 1.0,
       tphhl$I$Z = 1.0,
       tplz$OE$Z = 1.0,
       tphz$OE$Z = 1.0,
       tpzh$OE$Z = 1.0,
       tpzl$OE$Z = 1.0;

     // path delays
     (OE *> Z) = (0, 0, tplz$OE$Z, tpzh$OE$Z, tphz$OE$Z, tpzl$OE$Z);
     (I *> Z) = (tpllh$I$Z, tphhl$I$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_NT02D4 (Z, I, OE);
input  I ;
input  OE ;
output Z ;

   bufif0 (Z, I, OE);

   specify
     // delay parameters
     specparam
       tpllh$I$Z = 1.0,
       tphhl$I$Z = 1.0,
       tplz$OE$Z = 1.0,
       tphz$OE$Z = 1.0,
       tpzh$OE$Z = 1.0,
       tpzl$OE$Z = 1.0;

     // path delays
     (OE *> Z) = (0, 0, tplz$OE$Z, tpzh$OE$Z, tphz$OE$Z, tpzl$OE$Z);
     (I *> Z) = (tpllh$I$Z, tphhl$I$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_NT02D6 (Z, I, OE);
input  I ;
input  OE ;
output Z ;

   bufif0 (Z, I, OE);

   specify
     // delay parameters
     specparam
       tpllh$I$Z = 1.0,
       tphhl$I$Z = 1.0,
       tplz$OE$Z = 1.0,
       tphz$OE$Z = 1.0,
       tpzh$OE$Z = 1.0,
       tpzl$OE$Z = 1.0;

     // path delays
     (OE *> Z) = (0, 0, tplz$OE$Z, tpzh$OE$Z, tphz$OE$Z, tpzl$OE$Z);
     (I *> Z) = (tpllh$I$Z, tphhl$I$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OA01D2 (Z, A1, A2, B);
input  A1 ;
input  A2 ;
input  B ;
output Z ;

   or  (I0_out, A1, A2);
   and (Z, I0_out, B);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$B$Z = 1.0,
       tphhl$B$Z = 1.0,
       tpllh$B$Z$A1_EQ_1_AN_A2_EQ_1 = 1.0,
       tphhl$B$Z$A1_EQ_1_AN_A2_EQ_1 = 1.0,
       tpllh$B$Z$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tphhl$B$Z$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tpllh$B$Z$A1_EQ_1_AN_A2_EQ_0 = 1.0,
       tphhl$B$Z$A1_EQ_1_AN_A2_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1)
       (B *> Z) = (tpllh$B$Z$A1_EQ_1_AN_A2_EQ_1, tphhl$B$Z$A1_EQ_1_AN_A2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0)
       (B *> Z) = (tpllh$B$Z$A1_EQ_1_AN_A2_EQ_0, tphhl$B$Z$A1_EQ_1_AN_A2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1)
       (B *> Z) = (tpllh$B$Z$A1_EQ_0_AN_A2_EQ_1, tphhl$B$Z$A1_EQ_0_AN_A2_EQ_1);
     ifnone
       (B *> Z) = (tpllh$B$Z,tphhl$B$Z);

     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OA01D4 (Z, A1, A2, B);
input  A1 ;
input  A2 ;
input  B ;
output Z ;

   or  (I0_out, A1, A2);
   and (Z, I0_out, B);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$B$Z = 1.0,
       tphhl$B$Z = 1.0,
       tpllh$B$Z$A1_EQ_1_AN_A2_EQ_1 = 1.0,
       tphhl$B$Z$A1_EQ_1_AN_A2_EQ_1 = 1.0,
       tpllh$B$Z$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tphhl$B$Z$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tpllh$B$Z$A1_EQ_1_AN_A2_EQ_0 = 1.0,
       tphhl$B$Z$A1_EQ_1_AN_A2_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1)
       (B *> Z) = (tpllh$B$Z$A1_EQ_1_AN_A2_EQ_1, tphhl$B$Z$A1_EQ_1_AN_A2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0)
       (B *> Z) = (tpllh$B$Z$A1_EQ_1_AN_A2_EQ_0, tphhl$B$Z$A1_EQ_1_AN_A2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1)
       (B *> Z) = (tpllh$B$Z$A1_EQ_0_AN_A2_EQ_1, tphhl$B$Z$A1_EQ_0_AN_A2_EQ_1);
     ifnone
       (B *> Z) = (tpllh$B$Z,tphhl$B$Z);

     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OA02D2 (Z, A1, A2, B1, B2);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
output Z ;

   or  (I0_out, B1, B2);
   or  (I1_out, A1, A2);
   and (Z, I0_out, I1_out);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$B1$Z = 1.0,
       tphhl$B1$Z = 1.0,
       tpllh$B2$Z = 1.0,
       tphhl$B2$Z = 1.0,
       tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0);
     ifnone
       (B2 *> Z) = (tpllh$B2$Z,tphhl$B2$Z);

     if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0);
     ifnone
       (B1 *> Z) = (tpllh$B1$Z,tphhl$B1$Z);

     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     ifnone
       (A2 *> Z) = (tpllh$A2$Z,tphhl$A2$Z);

     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     ifnone
       (A1 *> Z) = (tpllh$A1$Z,tphhl$A1$Z);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OA02D4 (Z, A1, A2, B1, B2);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
output Z ;

   or  (I0_out, B1, B2);
   or  (I1_out, A1, A2);
   and (Z, I0_out, I1_out);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$B1$Z = 1.0,
       tphhl$B1$Z = 1.0,
       tpllh$B2$Z = 1.0,
       tphhl$B2$Z = 1.0,
       tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0);
     ifnone
       (B2 *> Z) = (tpllh$B2$Z,tphhl$B2$Z);

     if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0);
     ifnone
       (B1 *> Z) = (tpllh$B1$Z,tphhl$B1$Z);

     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     ifnone
       (A2 *> Z) = (tpllh$A2$Z,tphhl$A2$Z);

     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     ifnone
       (A1 *> Z) = (tpllh$A1$Z,tphhl$A1$Z);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OA03D2 (Z, A1, A2, A3, B);
input  A1 ;
input  A2 ;
input  A3 ;
input  B ;
output Z ;

   or  (I1_out, A1, A2, A3);
   and (Z, I1_out, B);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$A3$Z = 1.0,
       tphhl$A3$Z = 1.0,
       tpllh$B$Z = 1.0,
       tphhl$B$Z = 1.0,
       tpllh$B$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1 = 1.0,
       tphhl$B$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1 = 1.0,
       tpllh$B$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1 = 1.0,
       tphhl$B$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1 = 1.0,
       tpllh$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0 = 1.0,
       tphhl$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0 = 1.0,
       tpllh$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0 = 1.0,
       tphhl$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
       (B *> Z) = (tpllh$B$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1, tphhl$B$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
       (B *> Z) = (tpllh$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0, tphhl$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
       (B *> Z) = (tpllh$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0, tphhl$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
       (B *> Z) = (tpllh$B$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1, tphhl$B$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1);
     ifnone
       (B *> Z) = (tpllh$B$Z,tphhl$B$Z);

     (A3 *> Z) = (tpllh$A3$Z, tphhl$A3$Z);
     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OA03D4 (Z, A1, A2, A3, B);
input  A1 ;
input  A2 ;
input  A3 ;
input  B ;
output Z ;

   or  (I1_out, A1, A2, A3);
   and (Z, I1_out, B);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$A3$Z = 1.0,
       tphhl$A3$Z = 1.0,
       tpllh$B$Z = 1.0,
       tphhl$B$Z = 1.0,
       tpllh$B$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1 = 1.0,
       tphhl$B$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1 = 1.0,
       tpllh$B$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1 = 1.0,
       tphhl$B$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1 = 1.0,
       tpllh$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0 = 1.0,
       tphhl$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0 = 1.0,
       tpllh$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0 = 1.0,
       tphhl$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
       (B *> Z) = (tpllh$B$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1, tphhl$B$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
       (B *> Z) = (tpllh$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0, tphhl$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
       (B *> Z) = (tpllh$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0, tphhl$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
       (B *> Z) = (tpllh$B$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1, tphhl$B$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1);
     ifnone
       (B *> Z) = (tpllh$B$Z,tphhl$B$Z);

     (A3 *> Z) = (tpllh$A3$Z, tphhl$A3$Z);
     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OA04D2 (Z, A1, A2, A3, B1, B2);
input  A1 ;
input  A2 ;
input  A3 ;
input  B1 ;
input  B2 ;
output Z ;

   or  (I1_out, A1, A2, A3);
   or  (I2_out, B1, B2);
   and (Z, I1_out, I2_out);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$A3$Z = 1.0,
       tphhl$A3$Z = 1.0,
       tpllh$B1$Z = 1.0,
       tphhl$B1$Z = 1.0,
       tpllh$B2$Z = 1.0,
       tphhl$B2$Z = 1.0,
       tpllh$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tpllh$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tpllh$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_0 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0);
     ifnone
       (B2 *> Z) = (tpllh$B2$Z,tphhl$B2$Z);

     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_0, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_0, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_0, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_0, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_0);
     ifnone
       (B1 *> Z) = (tpllh$B1$Z,tphhl$B1$Z);

     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (A3 *> Z) = (tpllh$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tphhl$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A3 *> Z) = (tpllh$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A3 *> Z) = (tpllh$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     ifnone
       (A3 *> Z) = (tpllh$A3$Z,tphhl$A3$Z);

     if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tphhl$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     ifnone
       (A2 *> Z) = (tpllh$A2$Z,tphhl$A2$Z);

     if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tphhl$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     ifnone
       (A1 *> Z) = (tpllh$A1$Z,tphhl$A1$Z);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OA04D4 (Z, A1, A2, A3, B1, B2);
input  A1 ;
input  A2 ;
input  A3 ;
input  B1 ;
input  B2 ;
output Z ;

   or  (I1_out, A1, A2, A3);
   or  (I2_out, B1, B2);
   and (Z, I1_out, I2_out);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$A3$Z = 1.0,
       tphhl$A3$Z = 1.0,
       tpllh$B1$Z = 1.0,
       tphhl$B1$Z = 1.0,
       tpllh$B2$Z = 1.0,
       tphhl$B2$Z = 1.0,
       tpllh$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tpllh$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tpllh$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_0 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0);
     ifnone
       (B2 *> Z) = (tpllh$B2$Z,tphhl$B2$Z);

     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_0, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_0, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_0, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_0, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_0);
     ifnone
       (B1 *> Z) = (tpllh$B1$Z,tphhl$B1$Z);

     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (A3 *> Z) = (tpllh$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tphhl$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A3 *> Z) = (tpllh$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A3 *> Z) = (tpllh$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     ifnone
       (A3 *> Z) = (tpllh$A3$Z,tphhl$A3$Z);

     if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tphhl$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     ifnone
       (A2 *> Z) = (tpllh$A2$Z,tphhl$A2$Z);

     if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tphhl$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     ifnone
       (A1 *> Z) = (tpllh$A1$Z,tphhl$A1$Z);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OA05D2 (Z, A1, A2, A3, B1, B2, B3);
input  A1 ;
input  A2 ;
input  A3 ;
input  B1 ;
input  B2 ;
input  B3 ;
output Z ;

   or  (I1_out, A1, A2, A3);
   or  (I3_out, B1, B2, B3);
   and (Z, I1_out, I3_out);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$A3$Z = 1.0,
       tphhl$A3$Z = 1.0,
       tpllh$B1$Z = 1.0,
       tphhl$B1$Z = 1.0,
       tpllh$B2$Z = 1.0,
       tphhl$B2$Z = 1.0,
       tpllh$B3$Z = 1.0,
       tphhl$B3$Z = 1.0,
       tpllh$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tpllh$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tpllh$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tpllh$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tpllh$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tphhl$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tpllh$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphhl$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tpllh$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tphhl$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tpllh$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphhl$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B3_EQ_0 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B3_EQ_0 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0_AN_B3_EQ_0 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0_AN_B3_EQ_0 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0_AN_B3_EQ_0 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0_AN_B3_EQ_0 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B3_EQ_0 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B3_EQ_0 = 1.0,
       tpllh$B3$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$B3$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tpllh$B3$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$B3$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tpllh$B3$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$B3$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tpllh$B3$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$B3$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (B3 *> Z) = (tpllh$B3$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tphhl$B3$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
       (B3 *> Z) = (tpllh$B3$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0, tphhl$B3$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
       (B3 *> Z) = (tpllh$B3$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0, tphhl$B3$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (B3 *> Z) = (tpllh$B3$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tphhl$B3$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (B3 *> Z) = (tpllh$B3$Z,tphhl$B3$Z);

     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B3_EQ_0, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B3_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B3_EQ_0, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B3_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0_AN_B3_EQ_0, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0_AN_B3_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0_AN_B3_EQ_0, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0_AN_B3_EQ_0);
     ifnone
       (B2 *> Z) = (tpllh$B2$Z,tphhl$B2$Z);

     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0);
     ifnone
       (B1 *> Z) = (tpllh$B1$Z,tphhl$B1$Z);

     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
       (A3 *> Z) = (tpllh$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1, tphhl$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
       (A3 *> Z) = (tpllh$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0, tphhl$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
       (A3 *> Z) = (tpllh$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0, tphhl$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
       (A3 *> Z) = (tpllh$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1, tphhl$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1);
     ifnone
       (A3 *> Z) = (tpllh$A3$Z,tphhl$A3$Z);

     if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1, tphhl$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0, tphhl$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0);
     if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0, tphhl$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0);
     if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1, tphhl$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1);
     ifnone
       (A2 *> Z) = (tpllh$A2$Z,tphhl$A2$Z);

     if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1, tphhl$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0, tphhl$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0);
     if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0, tphhl$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0);
     if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1, tphhl$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1);
     ifnone
       (A1 *> Z) = (tpllh$A1$Z,tphhl$A1$Z);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OA05D4 (Z, A1, A2, A3, B1, B2, B3);
input  A1 ;
input  A2 ;
input  A3 ;
input  B1 ;
input  B2 ;
input  B3 ;
output Z ;

   or  (I1_out, A1, A2, A3);
   or  (I3_out, B1, B2, B3);
   and (Z, I1_out, I3_out);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$A3$Z = 1.0,
       tphhl$A3$Z = 1.0,
       tpllh$B1$Z = 1.0,
       tphhl$B1$Z = 1.0,
       tpllh$B2$Z = 1.0,
       tphhl$B2$Z = 1.0,
       tpllh$B3$Z = 1.0,
       tphhl$B3$Z = 1.0,
       tpllh$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tpllh$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tpllh$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tpllh$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tpllh$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tphhl$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tpllh$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphhl$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tpllh$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tphhl$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tpllh$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphhl$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B3_EQ_0 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B3_EQ_0 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0_AN_B3_EQ_0 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0_AN_B3_EQ_0 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0_AN_B3_EQ_0 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0_AN_B3_EQ_0 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B3_EQ_0 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B3_EQ_0 = 1.0,
       tpllh$B3$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$B3$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tpllh$B3$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$B3$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tpllh$B3$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$B3$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tpllh$B3$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$B3$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (B3 *> Z) = (tpllh$B3$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tphhl$B3$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
       (B3 *> Z) = (tpllh$B3$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0, tphhl$B3$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
       (B3 *> Z) = (tpllh$B3$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0, tphhl$B3$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (B3 *> Z) = (tpllh$B3$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tphhl$B3$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (B3 *> Z) = (tpllh$B3$Z,tphhl$B3$Z);

     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B3_EQ_0, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B3_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B3_EQ_0, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B3_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0_AN_B3_EQ_0, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0_AN_B3_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0_AN_B3_EQ_0, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0_AN_B3_EQ_0);
     ifnone
       (B2 *> Z) = (tpllh$B2$Z,tphhl$B2$Z);

     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0);
     ifnone
       (B1 *> Z) = (tpllh$B1$Z,tphhl$B1$Z);

     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
       (A3 *> Z) = (tpllh$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1, tphhl$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
       (A3 *> Z) = (tpllh$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0, tphhl$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
       (A3 *> Z) = (tpllh$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0, tphhl$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
       (A3 *> Z) = (tpllh$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1, tphhl$A3$Z$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1);
     ifnone
       (A3 *> Z) = (tpllh$A3$Z,tphhl$A3$Z);

     if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1, tphhl$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0, tphhl$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0);
     if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0, tphhl$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0);
     if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1, tphhl$A2$Z$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1);
     ifnone
       (A2 *> Z) = (tpllh$A2$Z,tphhl$A2$Z);

     if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1, tphhl$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0, tphhl$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0);
     if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0, tphhl$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0);
     if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1, tphhl$A1$Z$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1);
     ifnone
       (A1 *> Z) = (tpllh$A1$Z,tphhl$A1$Z);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OA06D2 (Z, A1, A2, B, C);
input  A1 ;
input  A2 ;
input  B ;
input  C ;
output Z ;

   or  (I0_out, A1, A2);
   and (Z, I0_out, B, C);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$B$Z = 1.0,
       tphhl$B$Z = 1.0,
       tpllh$C$Z = 1.0,
       tphhl$C$Z = 1.0,
       tpllh$B$Z$A1_EQ_1_AN_A2_EQ_1_AN_C_EQ_1 = 1.0,
       tphhl$B$Z$A1_EQ_1_AN_A2_EQ_1_AN_C_EQ_1 = 1.0,
       tpllh$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_1 = 1.0,
       tphhl$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_1 = 1.0,
       tpllh$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_1 = 1.0,
       tphhl$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_1 = 1.0,
       tpllh$C$Z$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_1 = 1.0,
       tphhl$C$Z$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_1 = 1.0,
       tpllh$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B_EQ_1 = 1.0,
       tphhl$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B_EQ_1 = 1.0,
       tpllh$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B_EQ_1 = 1.0,
       tphhl$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B_EQ_1 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && B == 1'b1)
       (C *> Z) = (tpllh$C$Z$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_1, tphhl$C$Z$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b1)
       (C *> Z) = (tpllh$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B_EQ_1, tphhl$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b1)
       (C *> Z) = (tpllh$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B_EQ_1, tphhl$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B_EQ_1);
     ifnone
       (C *> Z) = (tpllh$C$Z,tphhl$C$Z);

     if (A1 == 1'b1 && A2 == 1'b1 && C == 1'b1)
       (B *> Z) = (tpllh$B$Z$A1_EQ_1_AN_A2_EQ_1_AN_C_EQ_1, tphhl$B$Z$A1_EQ_1_AN_A2_EQ_1_AN_C_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b1)
       (B *> Z) = (tpllh$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_1, tphhl$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b1)
       (B *> Z) = (tpllh$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_1, tphhl$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_1);
     ifnone
       (B *> Z) = (tpllh$B$Z,tphhl$B$Z);

     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OA06D4 (Z, A1, A2, B, C);
input  A1 ;
input  A2 ;
input  B ;
input  C ;
output Z ;

   or  (I0_out, A1, A2);
   and (Z, I0_out, B, C);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$B$Z = 1.0,
       tphhl$B$Z = 1.0,
       tpllh$C$Z = 1.0,
       tphhl$C$Z = 1.0,
       tpllh$B$Z$A1_EQ_1_AN_A2_EQ_1_AN_C_EQ_1 = 1.0,
       tphhl$B$Z$A1_EQ_1_AN_A2_EQ_1_AN_C_EQ_1 = 1.0,
       tpllh$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_1 = 1.0,
       tphhl$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_1 = 1.0,
       tpllh$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_1 = 1.0,
       tphhl$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_1 = 1.0,
       tpllh$C$Z$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_1 = 1.0,
       tphhl$C$Z$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_1 = 1.0,
       tpllh$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B_EQ_1 = 1.0,
       tphhl$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B_EQ_1 = 1.0,
       tpllh$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B_EQ_1 = 1.0,
       tphhl$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B_EQ_1 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && B == 1'b1)
       (C *> Z) = (tpllh$C$Z$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_1, tphhl$C$Z$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b1)
       (C *> Z) = (tpllh$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B_EQ_1, tphhl$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b1)
       (C *> Z) = (tpllh$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B_EQ_1, tphhl$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B_EQ_1);
     ifnone
       (C *> Z) = (tpllh$C$Z,tphhl$C$Z);

     if (A1 == 1'b1 && A2 == 1'b1 && C == 1'b1)
       (B *> Z) = (tpllh$B$Z$A1_EQ_1_AN_A2_EQ_1_AN_C_EQ_1, tphhl$B$Z$A1_EQ_1_AN_A2_EQ_1_AN_C_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b1)
       (B *> Z) = (tpllh$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_1, tphhl$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b1)
       (B *> Z) = (tpllh$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_1, tphhl$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_1);
     ifnone
       (B *> Z) = (tpllh$B$Z,tphhl$B$Z);

     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OA07D2 (Z, A1, A2, B1, B2, C);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
input  C ;
output Z ;

   or  (I0_out, A1, A2);
   or  (I1_out, B1, B2);
   and (Z, I0_out, I1_out, C);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$B1$Z = 1.0,
       tphhl$B1$Z = 1.0,
       tpllh$B2$Z = 1.0,
       tphhl$B2$Z = 1.0,
       tpllh$C$Z = 1.0,
       tphhl$C$Z = 1.0,
       tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_1 = 1.0,
       tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C_EQ_1 = 1.0,
       tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_C_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_C_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C_EQ_1 = 1.0,
       tpllh$C$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$C$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tpllh$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
       (C *> Z) = (tpllh$C$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1, tphhl$C$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (C *> Z) = (tpllh$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (C *> Z) = (tpllh$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (C *> Z) = (tpllh$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (C *> Z) = (tpllh$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     ifnone
       (C *> Z) = (tpllh$C$Z,tphhl$C$Z);

     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_C_EQ_1, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_C_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C_EQ_1, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C_EQ_1, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C_EQ_1);
     ifnone
       (B2 *> Z) = (tpllh$B2$Z,tphhl$B2$Z);

     if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0_AN_C_EQ_1, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0_AN_C_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C_EQ_1, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C_EQ_1, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C_EQ_1);
     ifnone
       (B1 *> Z) = (tpllh$B1$Z,tphhl$B1$Z);

     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C_EQ_1, tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C_EQ_1);
     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_1, tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_1);
     if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_1, tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_1);
     ifnone
       (A2 *> Z) = (tpllh$A2$Z,tphhl$A2$Z);

     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C_EQ_1, tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C_EQ_1);
     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_1, tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_1);
     if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_1, tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_1);
     ifnone
       (A1 *> Z) = (tpllh$A1$Z,tphhl$A1$Z);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OA07D4 (Z, A1, A2, B1, B2, C);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
input  C ;
output Z ;

   or  (I0_out, A1, A2);
   or  (I1_out, B1, B2);
   and (Z, I0_out, I1_out, C);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$B1$Z = 1.0,
       tphhl$B1$Z = 1.0,
       tpllh$B2$Z = 1.0,
       tphhl$B2$Z = 1.0,
       tpllh$C$Z = 1.0,
       tphhl$C$Z = 1.0,
       tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_1 = 1.0,
       tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C_EQ_1 = 1.0,
       tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_C_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_C_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C_EQ_1 = 1.0,
       tpllh$C$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$C$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tpllh$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
       (C *> Z) = (tpllh$C$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1, tphhl$C$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (C *> Z) = (tpllh$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (C *> Z) = (tpllh$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$C$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (C *> Z) = (tpllh$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (C *> Z) = (tpllh$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$C$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     ifnone
       (C *> Z) = (tpllh$C$Z,tphhl$C$Z);

     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_C_EQ_1, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_C_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C_EQ_1, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C_EQ_1, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C_EQ_1);
     ifnone
       (B2 *> Z) = (tpllh$B2$Z,tphhl$B2$Z);

     if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0_AN_C_EQ_1, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0_AN_C_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C_EQ_1, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C_EQ_1, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C_EQ_1);
     ifnone
       (B1 *> Z) = (tpllh$B1$Z,tphhl$B1$Z);

     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C_EQ_1, tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C_EQ_1);
     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_1, tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_1);
     if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_1, tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_1);
     ifnone
       (A2 *> Z) = (tpllh$A2$Z,tphhl$A2$Z);

     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C_EQ_1, tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C_EQ_1);
     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_1, tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_1);
     if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_1, tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_1);
     ifnone
       (A1 *> Z) = (tpllh$A1$Z,tphhl$A1$Z);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OA08D2 (Z, A1, A2, B1, B2, C1, C2);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
input  C1 ;
input  C2 ;
output Z ;

   or  (I0_out, C1, C2);
   or  (I1_out, A1, A2);
   or  (I3_out, B1, B2);
   and (Z, I0_out, I1_out, I3_out);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$B1$Z = 1.0,
       tphhl$B1$Z = 1.0,
       tpllh$B2$Z = 1.0,
       tphhl$B2$Z = 1.0,
       tpllh$C1$Z = 1.0,
       tphhl$C1$Z = 1.0,
       tpllh$C2$Z = 1.0,
       tphhl$C2$Z = 1.0,
       tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_1 = 1.0,
       tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_1 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tpllh$C1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_C2_EQ_0 = 1.0,
       tphhl$C1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_C2_EQ_0 = 1.0,
       tpllh$C1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_0 = 1.0,
       tphhl$C1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_0 = 1.0,
       tpllh$C1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_0 = 1.0,
       tphhl$C1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_0 = 1.0,
       tpllh$C1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_0 = 1.0,
       tphhl$C1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_0 = 1.0,
       tpllh$C1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_0 = 1.0,
       tphhl$C1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_0 = 1.0,
       tpllh$C2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_0 = 1.0,
       tphhl$C2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_0 = 1.0,
       tpllh$C2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0 = 1.0,
       tphhl$C2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0 = 1.0,
       tpllh$C2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0 = 1.0,
       tphhl$C2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0 = 1.0,
       tpllh$C2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0 = 1.0,
       tphhl$C2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0 = 1.0,
       tpllh$C2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0 = 1.0,
       tphhl$C2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
       (C2 *> Z) = (tpllh$C2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_0, tphhl$C2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
       (C2 *> Z) = (tpllh$C2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0, tphhl$C2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
       (C2 *> Z) = (tpllh$C2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0, tphhl$C2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
       (C2 *> Z) = (tpllh$C2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0, tphhl$C2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
       (C2 *> Z) = (tpllh$C2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0, tphhl$C2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0);
     ifnone
       (C2 *> Z) = (tpllh$C2$Z,tphhl$C2$Z);

     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
       (C1 *> Z) = (tpllh$C1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_C2_EQ_0, tphhl$C1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
       (C1 *> Z) = (tpllh$C1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_0, tphhl$C1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
       (C1 *> Z) = (tpllh$C1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_0, tphhl$C1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
       (C1 *> Z) = (tpllh$C1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_0, tphhl$C1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
       (C1 *> Z) = (tpllh$C1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_0, tphhl$C1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_0);
     ifnone
       (C1 *> Z) = (tpllh$C1$Z,tphhl$C1$Z);

     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_1, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1);
     ifnone
       (B2 *> Z) = (tpllh$B2$Z,tphhl$B2$Z);

     if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_1, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1);
     ifnone
       (B1 *> Z) = (tpllh$B1$Z,tphhl$B1$Z);

     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_1, tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_1);
     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0, tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1, tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0, tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1, tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1);
     ifnone
       (A2 *> Z) = (tpllh$A2$Z,tphhl$A2$Z);

     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_1, tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_1);
     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0, tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1, tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0, tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1, tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1);
     ifnone
       (A1 *> Z) = (tpllh$A1$Z,tphhl$A1$Z);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OA08D4 (Z, A1, A2, B1, B2, C1, C2);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
input  C1 ;
input  C2 ;
output Z ;

   or  (I0_out, C1, C2);
   or  (I1_out, A1, A2);
   or  (I3_out, B1, B2);
   and (Z, I0_out, I1_out, I3_out);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$B1$Z = 1.0,
       tphhl$B1$Z = 1.0,
       tpllh$B2$Z = 1.0,
       tphhl$B2$Z = 1.0,
       tpllh$C1$Z = 1.0,
       tphhl$C1$Z = 1.0,
       tpllh$C2$Z = 1.0,
       tphhl$C2$Z = 1.0,
       tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_1 = 1.0,
       tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_1 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tpllh$C1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_C2_EQ_0 = 1.0,
       tphhl$C1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_C2_EQ_0 = 1.0,
       tpllh$C1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_0 = 1.0,
       tphhl$C1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_0 = 1.0,
       tpllh$C1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_0 = 1.0,
       tphhl$C1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_0 = 1.0,
       tpllh$C1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_0 = 1.0,
       tphhl$C1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_0 = 1.0,
       tpllh$C1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_0 = 1.0,
       tphhl$C1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_0 = 1.0,
       tpllh$C2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_0 = 1.0,
       tphhl$C2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_0 = 1.0,
       tpllh$C2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0 = 1.0,
       tphhl$C2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0 = 1.0,
       tpllh$C2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0 = 1.0,
       tphhl$C2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0 = 1.0,
       tpllh$C2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0 = 1.0,
       tphhl$C2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0 = 1.0,
       tpllh$C2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0 = 1.0,
       tphhl$C2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
       (C2 *> Z) = (tpllh$C2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_0, tphhl$C2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
       (C2 *> Z) = (tpllh$C2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0, tphhl$C2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
       (C2 *> Z) = (tpllh$C2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0, tphhl$C2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
       (C2 *> Z) = (tpllh$C2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0, tphhl$C2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
       (C2 *> Z) = (tpllh$C2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0, tphhl$C2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0);
     ifnone
       (C2 *> Z) = (tpllh$C2$Z,tphhl$C2$Z);

     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
       (C1 *> Z) = (tpllh$C1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_C2_EQ_0, tphhl$C1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
       (C1 *> Z) = (tpllh$C1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_0, tphhl$C1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
       (C1 *> Z) = (tpllh$C1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_0, tphhl$C1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
       (C1 *> Z) = (tpllh$C1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_0, tphhl$C1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
       (C1 *> Z) = (tpllh$C1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_0, tphhl$C1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_0);
     ifnone
       (C1 *> Z) = (tpllh$C1$Z,tphhl$C1$Z);

     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_1, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1, tphhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
       (B2 *> Z) = (tpllh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1, tphhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1);
     ifnone
       (B2 *> Z) = (tpllh$B2$Z,tphhl$B2$Z);

     if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_1, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1, tphhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
       (B1 *> Z) = (tpllh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1, tphhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1);
     ifnone
       (B1 *> Z) = (tpllh$B1$Z,tphhl$B1$Z);

     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_1, tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_1);
     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0, tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1, tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0, tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1, tphhl$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1);
     ifnone
       (A2 *> Z) = (tpllh$A2$Z,tphhl$A2$Z);

     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_1, tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_1);
     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0, tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1, tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0, tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1, tphhl$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1);
     ifnone
       (A1 *> Z) = (tpllh$A1$Z,tphhl$A1$Z);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OAN1BBD1 (ZN, A1N, A2N, B);
input  A1N ;
input  A2N ;
input  B ;
output ZN ;

   and (I0_out, A1N, A2N);
   not (I1_out, I0_out);
   and (I2_out, I1_out, B);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tpllh$A1N$ZN = 1.0,
       tphhl$A1N$ZN = 1.0,
       tpllh$A2N$ZN = 1.0,
       tphhl$A2N$ZN = 1.0,
       tplhl$B$ZN = 1.0,
       tphlh$B$ZN = 1.0,
       tplhl$B$ZN$A1N_EQ_0_AN_A2N_EQ_0 = 1.0,
       tphlh$B$ZN$A1N_EQ_0_AN_A2N_EQ_0 = 1.0,
       tplhl$B$ZN$A1N_EQ_1_AN_A2N_EQ_0 = 1.0,
       tphlh$B$ZN$A1N_EQ_1_AN_A2N_EQ_0 = 1.0,
       tplhl$B$ZN$A1N_EQ_0_AN_A2N_EQ_1 = 1.0,
       tphlh$B$ZN$A1N_EQ_0_AN_A2N_EQ_1 = 1.0;

     // path delays
     if (A1N == 1'b1 && A2N == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1N_EQ_1_AN_A2N_EQ_0, tplhl$B$ZN$A1N_EQ_1_AN_A2N_EQ_0);
     if (A1N == 1'b0 && A2N == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1N_EQ_0_AN_A2N_EQ_1, tplhl$B$ZN$A1N_EQ_0_AN_A2N_EQ_1);
     if (A1N == 1'b0 && A2N == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1N_EQ_0_AN_A2N_EQ_0, tplhl$B$ZN$A1N_EQ_0_AN_A2N_EQ_0);
     ifnone
       (B *> ZN) = (tphlh$B$ZN,tplhl$B$ZN);

     (A2N *> ZN) = (tpllh$A2N$ZN, tphhl$A2N$ZN);
     (A1N *> ZN) = (tpllh$A1N$ZN, tphhl$A1N$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OAN1BBD2 (ZN, A1N, A2N, B);
input  A1N ;
input  A2N ;
input  B ;
output ZN ;

   and (I0_out, A1N, A2N);
   not (I1_out, I0_out);
   and (I2_out, I1_out, B);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tpllh$A1N$ZN = 1.0,
       tphhl$A1N$ZN = 1.0,
       tpllh$A2N$ZN = 1.0,
       tphhl$A2N$ZN = 1.0,
       tplhl$B$ZN = 1.0,
       tphlh$B$ZN = 1.0,
       tplhl$B$ZN$A1N_EQ_0_AN_A2N_EQ_0 = 1.0,
       tphlh$B$ZN$A1N_EQ_0_AN_A2N_EQ_0 = 1.0,
       tplhl$B$ZN$A1N_EQ_1_AN_A2N_EQ_0 = 1.0,
       tphlh$B$ZN$A1N_EQ_1_AN_A2N_EQ_0 = 1.0,
       tplhl$B$ZN$A1N_EQ_0_AN_A2N_EQ_1 = 1.0,
       tphlh$B$ZN$A1N_EQ_0_AN_A2N_EQ_1 = 1.0;

     // path delays
     if (A1N == 1'b1 && A2N == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1N_EQ_1_AN_A2N_EQ_0, tplhl$B$ZN$A1N_EQ_1_AN_A2N_EQ_0);
     if (A1N == 1'b0 && A2N == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1N_EQ_0_AN_A2N_EQ_1, tplhl$B$ZN$A1N_EQ_0_AN_A2N_EQ_1);
     if (A1N == 1'b0 && A2N == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1N_EQ_0_AN_A2N_EQ_0, tplhl$B$ZN$A1N_EQ_0_AN_A2N_EQ_0);
     ifnone
       (B *> ZN) = (tphlh$B$ZN,tplhl$B$ZN);

     (A2N *> ZN) = (tpllh$A2N$ZN, tphhl$A2N$ZN);
     (A1N *> ZN) = (tpllh$A1N$ZN, tphhl$A1N$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OAN1BBD4 (ZN, A1N, A2N, B);
input  A1N ;
input  A2N ;
input  B ;
output ZN ;

   and (I0_out, A1N, A2N);
   not (I1_out, I0_out);
   and (I2_out, I1_out, B);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tpllh$A1N$ZN = 1.0,
       tphhl$A1N$ZN = 1.0,
       tpllh$A2N$ZN = 1.0,
       tphhl$A2N$ZN = 1.0,
       tplhl$B$ZN = 1.0,
       tphlh$B$ZN = 1.0,
       tplhl$B$ZN$A1N_EQ_0_AN_A2N_EQ_0 = 1.0,
       tphlh$B$ZN$A1N_EQ_0_AN_A2N_EQ_0 = 1.0,
       tplhl$B$ZN$A1N_EQ_1_AN_A2N_EQ_0 = 1.0,
       tphlh$B$ZN$A1N_EQ_1_AN_A2N_EQ_0 = 1.0,
       tplhl$B$ZN$A1N_EQ_0_AN_A2N_EQ_1 = 1.0,
       tphlh$B$ZN$A1N_EQ_0_AN_A2N_EQ_1 = 1.0;

     // path delays
     if (A1N == 1'b1 && A2N == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1N_EQ_1_AN_A2N_EQ_0, tplhl$B$ZN$A1N_EQ_1_AN_A2N_EQ_0);
     if (A1N == 1'b0 && A2N == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1N_EQ_0_AN_A2N_EQ_1, tplhl$B$ZN$A1N_EQ_0_AN_A2N_EQ_1);
     if (A1N == 1'b0 && A2N == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1N_EQ_0_AN_A2N_EQ_0, tplhl$B$ZN$A1N_EQ_0_AN_A2N_EQ_0);
     ifnone
       (B *> ZN) = (tphlh$B$ZN,tplhl$B$ZN);

     (A2N *> ZN) = (tpllh$A2N$ZN, tphhl$A2N$ZN);
     (A1N *> ZN) = (tpllh$A1N$ZN, tphhl$A1N$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OAN1BD1 (ZN, A1, A2, BN);
input  A1 ;
input  A2 ;
input  BN ;
output ZN ;

   or  (I0_out, A1, A2);
   not (I1_out, I0_out);
   or  (ZN, I1_out, BN);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tpllh$BN$ZN = 1.0,
       tphhl$BN$ZN = 1.0,
       tpllh$BN$ZN$A1_EQ_1_AN_A2_EQ_1 = 1.0,
       tphhl$BN$ZN$A1_EQ_1_AN_A2_EQ_1 = 1.0,
       tpllh$BN$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tphhl$BN$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tpllh$BN$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0,
       tphhl$BN$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1)
       (BN *> ZN) = (tpllh$BN$ZN$A1_EQ_1_AN_A2_EQ_1, tphhl$BN$ZN$A1_EQ_1_AN_A2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0)
       (BN *> ZN) = (tpllh$BN$ZN$A1_EQ_1_AN_A2_EQ_0, tphhl$BN$ZN$A1_EQ_1_AN_A2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1)
       (BN *> ZN) = (tpllh$BN$ZN$A1_EQ_0_AN_A2_EQ_1, tphhl$BN$ZN$A1_EQ_0_AN_A2_EQ_1);
     ifnone
       (BN *> ZN) = (tpllh$BN$ZN,tphhl$BN$ZN);

     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OAN1BD2 (ZN, A1, A2, BN);
input  A1 ;
input  A2 ;
input  BN ;
output ZN ;

   or  (I0_out, A1, A2);
   not (I1_out, I0_out);
   or  (ZN, I1_out, BN);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tpllh$BN$ZN = 1.0,
       tphhl$BN$ZN = 1.0,
       tpllh$BN$ZN$A1_EQ_1_AN_A2_EQ_1 = 1.0,
       tphhl$BN$ZN$A1_EQ_1_AN_A2_EQ_1 = 1.0,
       tpllh$BN$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tphhl$BN$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tpllh$BN$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0,
       tphhl$BN$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1)
       (BN *> ZN) = (tpllh$BN$ZN$A1_EQ_1_AN_A2_EQ_1, tphhl$BN$ZN$A1_EQ_1_AN_A2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0)
       (BN *> ZN) = (tpllh$BN$ZN$A1_EQ_1_AN_A2_EQ_0, tphhl$BN$ZN$A1_EQ_1_AN_A2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1)
       (BN *> ZN) = (tpllh$BN$ZN$A1_EQ_0_AN_A2_EQ_1, tphhl$BN$ZN$A1_EQ_0_AN_A2_EQ_1);
     ifnone
       (BN *> ZN) = (tpllh$BN$ZN,tphhl$BN$ZN);

     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OAN1BD4 (ZN, A1, A2, BN);
input  A1 ;
input  A2 ;
input  BN ;
output ZN ;

   or  (I0_out, A1, A2);
   not (I1_out, I0_out);
   or  (ZN, I1_out, BN);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tpllh$BN$ZN = 1.0,
       tphhl$BN$ZN = 1.0,
       tpllh$BN$ZN$A1_EQ_1_AN_A2_EQ_1 = 1.0,
       tphhl$BN$ZN$A1_EQ_1_AN_A2_EQ_1 = 1.0,
       tpllh$BN$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tphhl$BN$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tpllh$BN$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0,
       tphhl$BN$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1)
       (BN *> ZN) = (tpllh$BN$ZN$A1_EQ_1_AN_A2_EQ_1, tphhl$BN$ZN$A1_EQ_1_AN_A2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0)
       (BN *> ZN) = (tpllh$BN$ZN$A1_EQ_1_AN_A2_EQ_0, tphhl$BN$ZN$A1_EQ_1_AN_A2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1)
       (BN *> ZN) = (tpllh$BN$ZN$A1_EQ_0_AN_A2_EQ_1, tphhl$BN$ZN$A1_EQ_0_AN_A2_EQ_1);
     ifnone
       (BN *> ZN) = (tpllh$BN$ZN,tphhl$BN$ZN);

     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OAN1D1 (ZN, A1, A2, B);
input  A1 ;
input  A2 ;
input  B ;
output ZN ;

   or  (I0_out, A1, A2);
   and (I1_out, I0_out, B);
   not (ZN, I1_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$B$ZN = 1.0,
       tphlh$B$ZN = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_1 = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_1, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1);
     ifnone
       (B *> ZN) = (tphlh$B$ZN,tplhl$B$ZN);

     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OAN1D2 (ZN, A1, A2, B);
input  A1 ;
input  A2 ;
input  B ;
output ZN ;

   or  (I0_out, A1, A2);
   and (I1_out, I0_out, B);
   not (ZN, I1_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$B$ZN = 1.0,
       tphlh$B$ZN = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_1 = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_1, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1);
     ifnone
       (B *> ZN) = (tphlh$B$ZN,tplhl$B$ZN);

     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OAN1D4 (ZN, A1, A2, B);
input  A1 ;
input  A2 ;
input  B ;
output ZN ;

   or  (I0_out, A1, A2);
   and (I1_out, I0_out, B);
   not (ZN, I1_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$B$ZN = 1.0,
       tphlh$B$ZN = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_1 = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_1, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1);
     ifnone
       (B *> ZN) = (tphlh$B$ZN,tplhl$B$ZN);

     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OAN2BBD1 (ZN, A1N, A2N, B1, B2);
input  A1N ;
input  A2N ;
input  B1 ;
input  B2 ;
output ZN ;

   and (I0_out, A1N, A2N);
   not (I1_out, I0_out);
   or  (I2_out, B1, B2);
   and (I3_out, I1_out, I2_out);
   not (ZN, I3_out);

   specify
     // delay parameters
     specparam
       tpllh$A1N$ZN = 1.0,
       tphhl$A1N$ZN = 1.0,
       tpllh$A2N$ZN = 1.0,
       tphhl$A2N$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tpllh$A1N$ZN$A2N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$A1N$ZN$A2N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tpllh$A1N$ZN$A2N_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A1N$ZN$A2N_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A1N$ZN$A2N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A1N$ZN$A2N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$A2N$ZN$A1N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$A2N$ZN$A1N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tpllh$A2N$ZN$A1N_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A2N$ZN$A1N_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A2N$ZN$A1N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A2N$ZN$A1N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1N_EQ_0_AN_A2N_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1N_EQ_0_AN_A2N_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$B2$ZN$A1N_EQ_0_AN_A2N_EQ_0_AN_B1_EQ_0 = 1.0,
       tphlh$B2$ZN$A1N_EQ_0_AN_A2N_EQ_0_AN_B1_EQ_0 = 1.0,
       tplhl$B2$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B1_EQ_0 = 1.0,
       tphlh$B2$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B1_EQ_0 = 1.0,
       tplhl$B2$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B1_EQ_0 = 1.0,
       tphlh$B2$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B1_EQ_0 = 1.0;

     // path delays
     if (A1N == 1'b1 && A2N == 1'b0 && B1 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B1_EQ_0, tplhl$B2$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B1_EQ_0);
     if (A1N == 1'b0 && A2N == 1'b1 && B1 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B1_EQ_0, tplhl$B2$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B1_EQ_0);
     if (A1N == 1'b0 && A2N == 1'b0 && B1 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1N_EQ_0_AN_A2N_EQ_0_AN_B1_EQ_0, tplhl$B2$ZN$A1N_EQ_0_AN_A2N_EQ_0_AN_B1_EQ_0);
     ifnone
       (B2 *> ZN) = (tphlh$B2$ZN,tplhl$B2$ZN);

     if (A1N == 1'b1 && A2N == 1'b0 && B2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B2_EQ_0, tplhl$B1$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B2_EQ_0);
     if (A1N == 1'b0 && A2N == 1'b1 && B2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B2_EQ_0, tplhl$B1$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B2_EQ_0);
     if (A1N == 1'b0 && A2N == 1'b0 && B2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1N_EQ_0_AN_A2N_EQ_0_AN_B2_EQ_0, tplhl$B1$ZN$A1N_EQ_0_AN_A2N_EQ_0_AN_B2_EQ_0);
     ifnone
       (B1 *> ZN) = (tphlh$B1$ZN,tplhl$B1$ZN);

     if (A1N == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
       (A2N *> ZN) = (tpllh$A2N$ZN$A1N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1, tphhl$A2N$ZN$A1N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1N == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A2N *> ZN) = (tpllh$A2N$ZN$A1N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A2N$ZN$A1N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1N == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A2N *> ZN) = (tpllh$A2N$ZN$A1N_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A2N$ZN$A1N_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     ifnone
       (A2N *> ZN) = (tpllh$A2N$ZN,tphhl$A2N$ZN);

     if (A2N == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
       (A1N *> ZN) = (tpllh$A1N$ZN$A2N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1, tphhl$A1N$ZN$A2N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A2N == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A1N *> ZN) = (tpllh$A1N$ZN$A2N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A1N$ZN$A2N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A2N == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A1N *> ZN) = (tpllh$A1N$ZN$A2N_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A1N$ZN$A2N_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     ifnone
       (A1N *> ZN) = (tpllh$A1N$ZN,tphhl$A1N$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OAN2BBD2 (ZN, A1N, A2N, B1, B2);
input  A1N ;
input  A2N ;
input  B1 ;
input  B2 ;
output ZN ;

   and (I0_out, A1N, A2N);
   not (I1_out, I0_out);
   or  (I2_out, B1, B2);
   and (I3_out, I1_out, I2_out);
   not (ZN, I3_out);

   specify
     // delay parameters
     specparam
       tpllh$A1N$ZN = 1.0,
       tphhl$A1N$ZN = 1.0,
       tpllh$A2N$ZN = 1.0,
       tphhl$A2N$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tpllh$A1N$ZN$A2N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$A1N$ZN$A2N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tpllh$A1N$ZN$A2N_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A1N$ZN$A2N_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A1N$ZN$A2N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A1N$ZN$A2N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$A2N$ZN$A1N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$A2N$ZN$A1N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tpllh$A2N$ZN$A1N_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A2N$ZN$A1N_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A2N$ZN$A1N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A2N$ZN$A1N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1N_EQ_0_AN_A2N_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1N_EQ_0_AN_A2N_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B2$ZN$A1N_EQ_0_AN_A2N_EQ_0_AN_B1_EQ_0 = 1.0,
       tphlh$B2$ZN$A1N_EQ_0_AN_A2N_EQ_0_AN_B1_EQ_0 = 1.0,
       tplhl$B2$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B1_EQ_0 = 1.0,
       tphlh$B2$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B1_EQ_0 = 1.0,
       tplhl$B2$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B1_EQ_0 = 1.0,
       tphlh$B2$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B1_EQ_0 = 1.0;

     // path delays
     if (A1N == 1'b1 && A2N == 1'b0 && B1 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B1_EQ_0, tplhl$B2$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B1_EQ_0);
     if (A1N == 1'b0 && A2N == 1'b1 && B1 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B1_EQ_0, tplhl$B2$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B1_EQ_0);
     if (A1N == 1'b0 && A2N == 1'b0 && B1 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1N_EQ_0_AN_A2N_EQ_0_AN_B1_EQ_0, tplhl$B2$ZN$A1N_EQ_0_AN_A2N_EQ_0_AN_B1_EQ_0);
     ifnone
       (B2 *> ZN) = (tphlh$B2$ZN,tplhl$B2$ZN);

     if (A1N == 1'b1 && A2N == 1'b0 && B2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B2_EQ_0, tplhl$B1$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B2_EQ_0);
     if (A1N == 1'b0 && A2N == 1'b1 && B2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B2_EQ_0, tplhl$B1$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B2_EQ_0);
     if (A1N == 1'b0 && A2N == 1'b0 && B2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1N_EQ_0_AN_A2N_EQ_0_AN_B2_EQ_0, tplhl$B1$ZN$A1N_EQ_0_AN_A2N_EQ_0_AN_B2_EQ_0);
     ifnone
       (B1 *> ZN) = (tphlh$B1$ZN,tplhl$B1$ZN);

     if (A1N == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
       (A2N *> ZN) = (tpllh$A2N$ZN$A1N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1, tphhl$A2N$ZN$A1N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1N == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A2N *> ZN) = (tpllh$A2N$ZN$A1N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A2N$ZN$A1N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1N == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A2N *> ZN) = (tpllh$A2N$ZN$A1N_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A2N$ZN$A1N_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     ifnone
       (A2N *> ZN) = (tpllh$A2N$ZN,tphhl$A2N$ZN);

     if (A2N == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
       (A1N *> ZN) = (tpllh$A1N$ZN$A2N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1, tphhl$A1N$ZN$A2N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A2N == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A1N *> ZN) = (tpllh$A1N$ZN$A2N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A1N$ZN$A2N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A2N == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A1N *> ZN) = (tpllh$A1N$ZN$A2N_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A1N$ZN$A2N_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     ifnone
       (A1N *> ZN) = (tpllh$A1N$ZN,tphhl$A1N$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OAN2BBD4 (ZN, A1N, A2N, B1, B2);
input  A1N ;
input  A2N ;
input  B1 ;
input  B2 ;
output ZN ;

   and (I0_out, A1N, A2N);
   not (I1_out, I0_out);
   or  (I2_out, B1, B2);
   and (I3_out, I1_out, I2_out);
   not (ZN, I3_out);

   specify
     // delay parameters
     specparam
       tpllh$A1N$ZN = 1.0,
       tphhl$A1N$ZN = 1.0,
       tpllh$A2N$ZN = 1.0,
       tphhl$A2N$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tpllh$A1N$ZN$A2N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$A1N$ZN$A2N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tpllh$A1N$ZN$A2N_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A1N$ZN$A2N_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A1N$ZN$A2N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A1N$ZN$A2N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$A2N$ZN$A1N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$A2N$ZN$A1N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tpllh$A2N$ZN$A1N_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A2N$ZN$A1N_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A2N$ZN$A1N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A2N$ZN$A1N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1N_EQ_0_AN_A2N_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1N_EQ_0_AN_A2N_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B2$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B1_EQ_0 = 1.0,
       tphlh$B2$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B1_EQ_0 = 1.0,
       tplhl$B2$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B1_EQ_0 = 1.0,
       tphlh$B2$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B1_EQ_0 = 1.0,
       tplhl$B2$ZN$A1N_EQ_0_AN_A2N_EQ_0_AN_B1_EQ_0 = 1.0,
       tphlh$B2$ZN$A1N_EQ_0_AN_A2N_EQ_0_AN_B1_EQ_0 = 1.0;

     // path delays
     if (A1N == 1'b1 && A2N == 1'b0 && B1 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B1_EQ_0, tplhl$B2$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B1_EQ_0);
     if (A1N == 1'b0 && A2N == 1'b1 && B1 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B1_EQ_0, tplhl$B2$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B1_EQ_0);
     if (A1N == 1'b0 && A2N == 1'b0 && B1 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1N_EQ_0_AN_A2N_EQ_0_AN_B1_EQ_0, tplhl$B2$ZN$A1N_EQ_0_AN_A2N_EQ_0_AN_B1_EQ_0);
     ifnone
       (B2 *> ZN) = (tphlh$B2$ZN,tplhl$B2$ZN);

     if (A1N == 1'b1 && A2N == 1'b0 && B2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B2_EQ_0, tplhl$B1$ZN$A1N_EQ_1_AN_A2N_EQ_0_AN_B2_EQ_0);
     if (A1N == 1'b0 && A2N == 1'b1 && B2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B2_EQ_0, tplhl$B1$ZN$A1N_EQ_0_AN_A2N_EQ_1_AN_B2_EQ_0);
     if (A1N == 1'b0 && A2N == 1'b0 && B2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1N_EQ_0_AN_A2N_EQ_0_AN_B2_EQ_0, tplhl$B1$ZN$A1N_EQ_0_AN_A2N_EQ_0_AN_B2_EQ_0);
     ifnone
       (B1 *> ZN) = (tphlh$B1$ZN,tplhl$B1$ZN);

     if (A1N == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
       (A2N *> ZN) = (tpllh$A2N$ZN$A1N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1, tphhl$A2N$ZN$A1N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1N == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A2N *> ZN) = (tpllh$A2N$ZN$A1N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A2N$ZN$A1N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1N == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A2N *> ZN) = (tpllh$A2N$ZN$A1N_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A2N$ZN$A1N_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     ifnone
       (A2N *> ZN) = (tpllh$A2N$ZN,tphhl$A2N$ZN);

     if (A2N == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
       (A1N *> ZN) = (tpllh$A1N$ZN$A2N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1, tphhl$A1N$ZN$A2N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A2N == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (A1N *> ZN) = (tpllh$A1N$ZN$A2N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A1N$ZN$A2N_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A2N == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (A1N *> ZN) = (tpllh$A1N$ZN$A2N_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A1N$ZN$A2N_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     ifnone
       (A1N *> ZN) = (tpllh$A1N$ZN,tphhl$A1N$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OAN2D1 (ZN, A1, A2, B1, B2);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
output ZN ;

   or  (I0_out, A1, A2);
   or  (I1_out, B1, B2);
   and (I2_out, I0_out, I1_out);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0);
     ifnone
       (B2 *> ZN) = (tphlh$B2$ZN,tplhl$B2$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0);
     ifnone
       (B1 *> ZN) = (tphlh$B1$ZN,tplhl$B1$ZN);

     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     ifnone
       (A2 *> ZN) = (tphlh$A2$ZN,tplhl$A2$ZN);

     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     ifnone
       (A1 *> ZN) = (tphlh$A1$ZN,tplhl$A1$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OAN2D2 (ZN, A1, A2, B1, B2);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
output ZN ;

   or  (I0_out, B1, B2);
   or  (I1_out, A1, A2);
   and (I2_out, I0_out, I1_out);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0);
     ifnone
       (B2 *> ZN) = (tphlh$B2$ZN,tplhl$B2$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0);
     ifnone
       (B1 *> ZN) = (tphlh$B1$ZN,tplhl$B1$ZN);

     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     ifnone
       (A2 *> ZN) = (tphlh$A2$ZN,tplhl$A2$ZN);

     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     ifnone
       (A1 *> ZN) = (tphlh$A1$ZN,tplhl$A1$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OAN2D4 (ZN, A1, A2, B1, B2);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
output ZN ;

   or  (I0_out, B1, B2);
   or  (I1_out, A1, A2);
   and (I2_out, I0_out, I1_out);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0);
     ifnone
       (B2 *> ZN) = (tphlh$B2$ZN,tplhl$B2$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0);
     ifnone
       (B1 *> ZN) = (tphlh$B1$ZN,tplhl$B1$ZN);

     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     ifnone
       (A2 *> ZN) = (tphlh$A2$ZN,tplhl$A2$ZN);

     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     ifnone
       (A1 *> ZN) = (tphlh$A1$ZN,tplhl$A1$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OAN3D1 (ZN, A1, A2, A3, B);
input  A1 ;
input  A2 ;
input  A3 ;
input  B ;
output ZN ;

   or  (I1_out, A1, A2, A3);
   and (I2_out, I1_out, B);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0,
       tplhl$B$ZN = 1.0,
       tphlh$B$ZN = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1 = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1 = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0 = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1);
     ifnone
       (B *> ZN) = (tphlh$B$ZN,tplhl$B$ZN);

     (A3 *> ZN) = (tphlh$A3$ZN, tplhl$A3$ZN);
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OAN3D2 (ZN, A1, A2, A3, B);
input  A1 ;
input  A2 ;
input  A3 ;
input  B ;
output ZN ;

   or  (I1_out, A1, A2, A3);
   and (I2_out, I1_out, B);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0,
       tplhl$B$ZN = 1.0,
       tphlh$B$ZN = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1 = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1 = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0 = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1);
     ifnone
       (B *> ZN) = (tphlh$B$ZN,tplhl$B$ZN);

     (A3 *> ZN) = (tphlh$A3$ZN, tplhl$A3$ZN);
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OAN3D4 (ZN, A1, A2, A3, B);
input  A1 ;
input  A2 ;
input  A3 ;
input  B ;
output ZN ;

   or  (I1_out, A1, A2, A3);
   and (I2_out, I1_out, B);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0,
       tplhl$B$ZN = 1.0,
       tphlh$B$ZN = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1 = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1 = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0 = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1);
     ifnone
       (B *> ZN) = (tphlh$B$ZN,tplhl$B$ZN);

     (A3 *> ZN) = (tphlh$A3$ZN, tplhl$A3$ZN);
     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OAN4D1 (ZN, A1, A2, A3, B1, B2);
input  A1 ;
input  A2 ;
input  A3 ;
input  B1 ;
input  B2 ;
output ZN ;

   or  (I0_out, B1, B2);
   or  (I2_out, A1, A2, A3);
   and (I3_out, I0_out, I2_out);
   not (ZN, I3_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0);
     ifnone
       (B2 *> ZN) = (tphlh$B2$ZN,tplhl$B2$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_0, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_0, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_0, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_0, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_0);
     ifnone
       (B1 *> ZN) = (tphlh$B1$ZN,tplhl$B1$ZN);

     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     ifnone
       (A3 *> ZN) = (tphlh$A3$ZN,tplhl$A3$ZN);

     if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     ifnone
       (A2 *> ZN) = (tphlh$A2$ZN,tplhl$A2$ZN);

     if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     ifnone
       (A1 *> ZN) = (tphlh$A1$ZN,tplhl$A1$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OAN4D2 (ZN, A1, A2, A3, B1, B2);
input  A1 ;
input  A2 ;
input  A3 ;
input  B1 ;
input  B2 ;
output ZN ;

   or  (I1_out, A1, A2, A3);
   or  (I2_out, B1, B2);
   and (I3_out, I1_out, I2_out);
   not (ZN, I3_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0);
     ifnone
       (B2 *> ZN) = (tphlh$B2$ZN,tplhl$B2$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_0, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_0, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_0, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_0, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_0);
     ifnone
       (B1 *> ZN) = (tphlh$B1$ZN,tplhl$B1$ZN);

     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     ifnone
       (A3 *> ZN) = (tphlh$A3$ZN,tplhl$A3$ZN);

     if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     ifnone
       (A2 *> ZN) = (tphlh$A2$ZN,tplhl$A2$ZN);

     if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     ifnone
       (A1 *> ZN) = (tphlh$A1$ZN,tplhl$A1$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OAN4D4 (ZN, A1, A2, A3, B1, B2);
input  A1 ;
input  A2 ;
input  A3 ;
input  B1 ;
input  B2 ;
output ZN ;

   or  (I1_out, A1, A2, A3);
   or  (I2_out, B1, B2);
   and (I3_out, I1_out, I2_out);
   not (ZN, I3_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0);
     ifnone
       (B2 *> ZN) = (tphlh$B2$ZN,tplhl$B2$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_0, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_0, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_0, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_0, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_0);
     ifnone
       (B1 *> ZN) = (tphlh$B1$ZN,tplhl$B1$ZN);

     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     ifnone
       (A3 *> ZN) = (tphlh$A3$ZN,tplhl$A3$ZN);

     if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     ifnone
       (A2 *> ZN) = (tphlh$A2$ZN,tplhl$A2$ZN);

     if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     ifnone
       (A1 *> ZN) = (tphlh$A1$ZN,tplhl$A1$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OAN5D1 (ZN, A1, A2, A3, B1, B2, B3);
input  A1 ;
input  A2 ;
input  A3 ;
input  B1 ;
input  B2 ;
input  B3 ;
output ZN ;

   or  (I1_out, B1, B2, B3);
   or  (I3_out, A1, A2, A3);
   and (I4_out, I1_out, I3_out);
   not (ZN, I4_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tplhl$B3$ZN = 1.0,
       tphlh$B3$ZN = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$B3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$B3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$B3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$B3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$B3$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$B3$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$B3$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$B3$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (B3 *> ZN) = (tphlh$B3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tplhl$B3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
       (B3 *> ZN) = (tphlh$B3$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0, tplhl$B3$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
       (B3 *> ZN) = (tphlh$B3$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0, tplhl$B3$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (B3 *> ZN) = (tphlh$B3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tplhl$B3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (B3 *> ZN) = (tphlh$B3$ZN,tplhl$B3$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B3_EQ_0, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B3_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B3_EQ_0, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B3_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0_AN_B3_EQ_0, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0_AN_B3_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0_AN_B3_EQ_0, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0_AN_B3_EQ_0);
     ifnone
       (B2 *> ZN) = (tphlh$B2$ZN,tplhl$B2$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0);
     ifnone
       (B1 *> ZN) = (tphlh$B1$ZN,tplhl$B1$ZN);

     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1, tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0, tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0, tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1, tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1);
     ifnone
       (A3 *> ZN) = (tphlh$A3$ZN,tplhl$A3$ZN);

     if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1, tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0, tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0);
     if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0, tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0);
     if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1, tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1);
     ifnone
       (A2 *> ZN) = (tphlh$A2$ZN,tplhl$A2$ZN);

     if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1, tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0, tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0);
     if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0, tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0);
     if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1, tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1);
     ifnone
       (A1 *> ZN) = (tphlh$A1$ZN,tplhl$A1$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OAN5D2 (ZN, A1, A2, A3, B1, B2, B3);
input  A1 ;
input  A2 ;
input  A3 ;
input  B1 ;
input  B2 ;
input  B3 ;
output ZN ;

   or  (I1_out, A1, A2, A3);
   or  (I3_out, B1, B2, B3);
   and (I4_out, I1_out, I3_out);
   not (ZN, I4_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tplhl$B3$ZN = 1.0,
       tphlh$B3$ZN = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$B3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$B3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$B3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$B3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$B3$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$B3$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$B3$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$B3$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (B3 *> ZN) = (tphlh$B3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tplhl$B3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
       (B3 *> ZN) = (tphlh$B3$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0, tplhl$B3$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
       (B3 *> ZN) = (tphlh$B3$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0, tplhl$B3$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (B3 *> ZN) = (tphlh$B3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tplhl$B3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (B3 *> ZN) = (tphlh$B3$ZN,tplhl$B3$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B3_EQ_0, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B3_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B3_EQ_0, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B3_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0_AN_B3_EQ_0, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0_AN_B3_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0_AN_B3_EQ_0, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0_AN_B3_EQ_0);
     ifnone
       (B2 *> ZN) = (tphlh$B2$ZN,tplhl$B2$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0);
     ifnone
       (B1 *> ZN) = (tphlh$B1$ZN,tplhl$B1$ZN);

     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1, tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0, tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0, tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1, tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1);
     ifnone
       (A3 *> ZN) = (tphlh$A3$ZN,tplhl$A3$ZN);

     if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1, tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0, tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0);
     if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0, tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0);
     if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1, tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1);
     ifnone
       (A2 *> ZN) = (tphlh$A2$ZN,tplhl$A2$ZN);

     if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1, tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0, tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0);
     if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0, tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0);
     if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1, tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1);
     ifnone
       (A1 *> ZN) = (tphlh$A1$ZN,tplhl$A1$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OAN5D4 (ZN, A1, A2, A3, B1, B2, B3);
input  A1 ;
input  A2 ;
input  A3 ;
input  B1 ;
input  B2 ;
input  B3 ;
output ZN ;

   or  (I1_out, A1, A2, A3);
   or  (I3_out, B1, B2, B3);
   and (I4_out, I1_out, I3_out);
   not (ZN, I4_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tplhl$B3$ZN = 1.0,
       tphlh$B3$ZN = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1 = 1.0,
       tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1 = 1.0,
       tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0 = 1.0,
       tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B3_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B3_EQ_0 = 1.0,
       tplhl$B3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$B3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$B3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$B3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$B3$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$B3$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$B3$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$B3$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (B3 *> ZN) = (tphlh$B3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tplhl$B3$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
       (B3 *> ZN) = (tphlh$B3$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0, tplhl$B3$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
       (B3 *> ZN) = (tphlh$B3$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0, tplhl$B3$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
       (B3 *> ZN) = (tphlh$B3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0, tplhl$B3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0_AN_B2_EQ_0);
     ifnone
       (B3 *> ZN) = (tphlh$B3$ZN,tplhl$B3$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B3_EQ_0, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B1_EQ_0_AN_B3_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B3_EQ_0, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B3_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0_AN_B3_EQ_0, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B1_EQ_0_AN_B3_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0_AN_B3_EQ_0, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B1_EQ_0_AN_B3_EQ_0);
     ifnone
       (B2 *> ZN) = (tphlh$B2$ZN,tplhl$B2$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_A3_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_A3_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_A3_EQ_0_AN_B2_EQ_0_AN_B3_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_0_AN_A3_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0);
     ifnone
       (B1 *> ZN) = (tphlh$B1$ZN,tplhl$B1$ZN);

     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1, tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0, tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0, tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1, tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1);
     ifnone
       (A3 *> ZN) = (tphlh$A3$ZN,tplhl$A3$ZN);

     if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1, tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0, tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0);
     if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0, tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0);
     if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1, tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1);
     ifnone
       (A2 *> ZN) = (tphlh$A2$ZN,tplhl$A2$ZN);

     if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1, tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_B3_EQ_1);
     if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0, tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_B3_EQ_0);
     if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0, tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_B3_EQ_0);
     if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1, tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0_AN_B1_EQ_0_AN_B2_EQ_0_AN_B3_EQ_1);
     ifnone
       (A1 *> ZN) = (tphlh$A1$ZN,tplhl$A1$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OAN6D1 (ZN, A1, A2, B, C);
input  A1 ;
input  A2 ;
input  B ;
input  C ;
output ZN ;

   or  (I0_out, A1, A2);
   and (I2_out, I0_out, B, C);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$B$ZN = 1.0,
       tphlh$B$ZN = 1.0,
       tplhl$C$ZN = 1.0,
       tphlh$C$ZN = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_C_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_C_EQ_1 = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_1 = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_1 = 1.0,
       tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_1 = 1.0,
       tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_1 = 1.0,
       tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B_EQ_1 = 1.0,
       tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B_EQ_1 = 1.0,
       tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B_EQ_1 = 1.0,
       tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B_EQ_1 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && B == 1'b1)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_1, tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b1)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B_EQ_1, tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b1)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B_EQ_1, tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B_EQ_1);
     ifnone
       (C *> ZN) = (tphlh$C$ZN,tplhl$C$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && C == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_C_EQ_1, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_C_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_1, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_1, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_1);
     ifnone
       (B *> ZN) = (tphlh$B$ZN,tplhl$B$ZN);

     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OAN6D2 (ZN, A1, A2, B, C);
input  A1 ;
input  A2 ;
input  B ;
input  C ;
output ZN ;

   or  (I0_out, A1, A2);
   and (I2_out, I0_out, B, C);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$B$ZN = 1.0,
       tphlh$B$ZN = 1.0,
       tplhl$C$ZN = 1.0,
       tphlh$C$ZN = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_C_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_C_EQ_1 = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_1 = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_1 = 1.0,
       tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_1 = 1.0,
       tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_1 = 1.0,
       tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B_EQ_1 = 1.0,
       tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B_EQ_1 = 1.0,
       tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B_EQ_1 = 1.0,
       tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B_EQ_1 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && B == 1'b1)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_1, tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b1)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B_EQ_1, tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b1)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B_EQ_1, tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B_EQ_1);
     ifnone
       (C *> ZN) = (tphlh$C$ZN,tplhl$C$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && C == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_C_EQ_1, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_C_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_1, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_1, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_1);
     ifnone
       (B *> ZN) = (tphlh$B$ZN,tplhl$B$ZN);

     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OAN6D4 (ZN, A1, A2, B, C);
input  A1 ;
input  A2 ;
input  B ;
input  C ;
output ZN ;

   or  (I0_out, A1, A2);
   and (I2_out, I0_out, B, C);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$B$ZN = 1.0,
       tphlh$B$ZN = 1.0,
       tplhl$C$ZN = 1.0,
       tphlh$C$ZN = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_C_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_C_EQ_1 = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_1 = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_1 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_1 = 1.0,
       tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_1 = 1.0,
       tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_1 = 1.0,
       tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B_EQ_1 = 1.0,
       tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B_EQ_1 = 1.0,
       tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B_EQ_1 = 1.0,
       tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B_EQ_1 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && B == 1'b1)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_1, tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b1)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B_EQ_1, tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b1)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B_EQ_1, tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B_EQ_1);
     ifnone
       (C *> ZN) = (tphlh$C$ZN,tplhl$C$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && C == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_C_EQ_1, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_C_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_1, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b1)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_1, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_1);
     ifnone
       (B *> ZN) = (tphlh$B$ZN,tplhl$B$ZN);

     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OAN7D1 (ZN, A1, A2, B1, B2, C);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
input  C ;
output ZN ;

   or  (I0_out, A1, A2);
   or  (I1_out, B1, B2);
   and (I3_out, I0_out, I1_out, C);
   not (ZN, I3_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tplhl$C$ZN = 1.0,
       tphlh$C$ZN = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_C_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_C_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C_EQ_1 = 1.0,
       tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1, tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     ifnone
       (C *> ZN) = (tphlh$C$ZN,tplhl$C$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_C_EQ_1, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_C_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C_EQ_1, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C_EQ_1, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C_EQ_1);
     ifnone
       (B2 *> ZN) = (tphlh$B2$ZN,tplhl$B2$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0_AN_C_EQ_1, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0_AN_C_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C_EQ_1, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C_EQ_1, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C_EQ_1);
     ifnone
       (B1 *> ZN) = (tphlh$B1$ZN,tplhl$B1$ZN);

     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C_EQ_1, tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C_EQ_1);
     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_1, tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_1);
     if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_1, tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_1);
     ifnone
       (A2 *> ZN) = (tphlh$A2$ZN,tplhl$A2$ZN);

     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C_EQ_1, tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C_EQ_1);
     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_1, tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_1);
     if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_1, tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_1);
     ifnone
       (A1 *> ZN) = (tphlh$A1$ZN,tplhl$A1$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OAN7D2 (ZN, A1, A2, B1, B2, C);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
input  C ;
output ZN ;

   or  (I0_out, A1, A2);
   or  (I1_out, B1, B2);
   and (I3_out, I0_out, I1_out, C);
   not (ZN, I3_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tplhl$C$ZN = 1.0,
       tphlh$C$ZN = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_C_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_C_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C_EQ_1 = 1.0,
       tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1, tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     ifnone
       (C *> ZN) = (tphlh$C$ZN,tplhl$C$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_C_EQ_1, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_C_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C_EQ_1, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C_EQ_1, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C_EQ_1);
     ifnone
       (B2 *> ZN) = (tphlh$B2$ZN,tplhl$B2$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0_AN_C_EQ_1, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0_AN_C_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C_EQ_1, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C_EQ_1, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C_EQ_1);
     ifnone
       (B1 *> ZN) = (tphlh$B1$ZN,tplhl$B1$ZN);

     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C_EQ_1, tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C_EQ_1);
     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_1, tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_1);
     if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_1, tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_1);
     ifnone
       (A2 *> ZN) = (tphlh$A2$ZN,tplhl$A2$ZN);

     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C_EQ_1, tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C_EQ_1);
     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_1, tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_1);
     if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_1, tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_1);
     ifnone
       (A1 *> ZN) = (tphlh$A1$ZN,tplhl$A1$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OAN7D4 (ZN, A1, A2, B1, B2, C);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
input  C ;
output ZN ;

   or  (I0_out, A1, A2);
   or  (I1_out, B1, B2);
   and (I3_out, I0_out, I1_out, C);
   not (ZN, I3_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tplhl$C$ZN = 1.0,
       tphlh$C$ZN = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_C_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_C_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C_EQ_1 = 1.0,
       tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1, tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1);
     ifnone
       (C *> ZN) = (tphlh$C$ZN,tplhl$C$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_C_EQ_1, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_C_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C_EQ_1, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C_EQ_1, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C_EQ_1);
     ifnone
       (B2 *> ZN) = (tphlh$B2$ZN,tplhl$B2$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0_AN_C_EQ_1, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0_AN_C_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C_EQ_1, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C_EQ_1, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C_EQ_1);
     ifnone
       (B1 *> ZN) = (tphlh$B1$ZN,tplhl$B1$ZN);

     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C_EQ_1, tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C_EQ_1);
     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_1, tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_1);
     if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_1, tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_1);
     ifnone
       (A2 *> ZN) = (tphlh$A2$ZN,tplhl$A2$ZN);

     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C_EQ_1, tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C_EQ_1);
     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_1, tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C_EQ_1);
     if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_1, tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C_EQ_1);
     ifnone
       (A1 *> ZN) = (tphlh$A1$ZN,tplhl$A1$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OAN8D1 (ZN, A1, A2, B1, B2, C1, C2);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
input  C1 ;
input  C2 ;
output ZN ;

   or  (I0_out, A1, A2);
   or  (I1_out, C1, C2);
   or  (I3_out, B1, B2);
   and (I4_out, I0_out, I1_out, I3_out);
   not (ZN, I4_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tplhl$C1$ZN = 1.0,
       tphlh$C1$ZN = 1.0,
       tplhl$C2$ZN = 1.0,
       tphlh$C2$ZN = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$C1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$C1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_0 = 1.0,
       tphlh$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_0 = 1.0,
       tplhl$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_0 = 1.0,
       tphlh$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_0 = 1.0,
       tplhl$C2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_0 = 1.0,
       tphlh$C2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_0 = 1.0,
       tplhl$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0 = 1.0,
       tphlh$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0 = 1.0,
       tplhl$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0 = 1.0,
       tphlh$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0 = 1.0,
       tplhl$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0 = 1.0,
       tphlh$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0 = 1.0,
       tplhl$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0 = 1.0,
       tphlh$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
       (C2 *> ZN) = (tphlh$C2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_0, tplhl$C2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
       (C2 *> ZN) = (tphlh$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0, tplhl$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
       (C2 *> ZN) = (tphlh$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0, tplhl$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
       (C2 *> ZN) = (tphlh$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0, tplhl$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
       (C2 *> ZN) = (tphlh$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0, tplhl$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0);
     ifnone
       (C2 *> ZN) = (tphlh$C2$ZN,tplhl$C2$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
       (C1 *> ZN) = (tphlh$C1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_C2_EQ_0, tplhl$C1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
       (C1 *> ZN) = (tphlh$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_0, tplhl$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
       (C1 *> ZN) = (tphlh$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_0, tplhl$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
       (C1 *> ZN) = (tphlh$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_0, tplhl$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
       (C1 *> ZN) = (tphlh$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_0, tplhl$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_0);
     ifnone
       (C1 *> ZN) = (tphlh$C1$ZN,tplhl$C1$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_1, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1);
     ifnone
       (B2 *> ZN) = (tphlh$B2$ZN,tplhl$B2$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_1, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1);
     ifnone
       (B1 *> ZN) = (tphlh$B1$ZN,tplhl$B1$ZN);

     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_1, tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_1);
     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1);
     ifnone
       (A2 *> ZN) = (tphlh$A2$ZN,tplhl$A2$ZN);

     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_1, tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_1);
     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1);
     ifnone
       (A1 *> ZN) = (tphlh$A1$ZN,tplhl$A1$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OAN8D2 (ZN, A1, A2, B1, B2, C1, C2);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
input  C1 ;
input  C2 ;
output ZN ;

   or  (I0_out, A1, A2);
   or  (I1_out, C1, C2);
   or  (I3_out, B1, B2);
   and (I4_out, I0_out, I1_out, I3_out);
   not (ZN, I4_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tplhl$C1$ZN = 1.0,
       tphlh$C1$ZN = 1.0,
       tplhl$C2$ZN = 1.0,
       tphlh$C2$ZN = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$C1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$C1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_0 = 1.0,
       tphlh$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_0 = 1.0,
       tplhl$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_0 = 1.0,
       tphlh$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_0 = 1.0,
       tplhl$C2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_0 = 1.0,
       tphlh$C2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_0 = 1.0,
       tplhl$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0 = 1.0,
       tphlh$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0 = 1.0,
       tplhl$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0 = 1.0,
       tphlh$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0 = 1.0,
       tplhl$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0 = 1.0,
       tphlh$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0 = 1.0,
       tplhl$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0 = 1.0,
       tphlh$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
       (C2 *> ZN) = (tphlh$C2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_0, tplhl$C2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
       (C2 *> ZN) = (tphlh$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0, tplhl$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
       (C2 *> ZN) = (tphlh$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0, tplhl$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
       (C2 *> ZN) = (tphlh$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0, tplhl$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
       (C2 *> ZN) = (tphlh$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0, tplhl$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0);
     ifnone
       (C2 *> ZN) = (tphlh$C2$ZN,tplhl$C2$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
       (C1 *> ZN) = (tphlh$C1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_C2_EQ_0, tplhl$C1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
       (C1 *> ZN) = (tphlh$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_0, tplhl$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
       (C1 *> ZN) = (tphlh$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_0, tplhl$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
       (C1 *> ZN) = (tphlh$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_0, tplhl$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
       (C1 *> ZN) = (tphlh$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_0, tplhl$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_0);
     ifnone
       (C1 *> ZN) = (tphlh$C1$ZN,tplhl$C1$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_1, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1);
     ifnone
       (B2 *> ZN) = (tphlh$B2$ZN,tplhl$B2$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_1, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1);
     ifnone
       (B1 *> ZN) = (tphlh$B1$ZN,tplhl$B1$ZN);

     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_1, tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_1);
     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1);
     ifnone
       (A2 *> ZN) = (tphlh$A2$ZN,tplhl$A2$ZN);

     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_1, tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_1);
     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1);
     ifnone
       (A1 *> ZN) = (tphlh$A1$ZN,tplhl$A1$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OAN8D4 (ZN, A1, A2, B1, B2, C1, C2);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
input  C1 ;
input  C2 ;
output ZN ;

   or  (I0_out, A1, A2);
   or  (I1_out, C1, C2);
   or  (I3_out, B1, B2);
   and (I4_out, I0_out, I1_out, I3_out);
   not (ZN, I4_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tplhl$C1$ZN = 1.0,
       tphlh$C1$ZN = 1.0,
       tplhl$C2$ZN = 1.0,
       tphlh$C2$ZN = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1 = 1.0,
       tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$C1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$C1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_0 = 1.0,
       tphlh$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_0 = 1.0,
       tplhl$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_0 = 1.0,
       tphlh$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_0 = 1.0,
       tplhl$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_0 = 1.0,
       tphlh$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_0 = 1.0,
       tplhl$C2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_0 = 1.0,
       tphlh$C2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_0 = 1.0,
       tplhl$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0 = 1.0,
       tphlh$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0 = 1.0,
       tplhl$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0 = 1.0,
       tphlh$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0 = 1.0,
       tplhl$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0 = 1.0,
       tphlh$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0 = 1.0,
       tplhl$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0 = 1.0,
       tphlh$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
       (C2 *> ZN) = (tphlh$C2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_0, tplhl$C2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
       (C2 *> ZN) = (tphlh$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0, tplhl$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
       (C2 *> ZN) = (tphlh$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0, tplhl$C2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
       (C2 *> ZN) = (tphlh$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0, tplhl$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
       (C2 *> ZN) = (tphlh$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0, tplhl$C2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0);
     ifnone
       (C2 *> ZN) = (tphlh$C2$ZN,tplhl$C2$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
       (C1 *> ZN) = (tphlh$C1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_C2_EQ_0, tplhl$C1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
       (C1 *> ZN) = (tphlh$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_0, tplhl$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
       (C1 *> ZN) = (tphlh$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_0, tplhl$C1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
       (C1 *> ZN) = (tphlh$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_0, tplhl$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_1_AN_B2_EQ_0_AN_C2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
       (C1 *> ZN) = (tphlh$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_0, tplhl$C1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_B2_EQ_1_AN_C2_EQ_0);
     ifnone
       (C1 *> ZN) = (tphlh$C1$ZN,tplhl$C1$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_1, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
       (B2 *> ZN) = (tphlh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1);
     ifnone
       (B2 *> ZN) = (tphlh$B2$ZN,tplhl$B2$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_1, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
       (B1 *> ZN) = (tphlh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1);
     ifnone
       (B1 *> ZN) = (tphlh$B1$ZN,tplhl$B1$ZN);

     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_1, tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_1);
     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1);
     ifnone
       (A2 *> ZN) = (tphlh$A2$ZN,tplhl$A2$ZN);

     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_1, tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_1);
     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0_AN_C1_EQ_0_AN_C2_EQ_1);
     if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0, tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_1_AN_C2_EQ_0);
     if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1, tplhl$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1_AN_C1_EQ_0_AN_C2_EQ_1);
     ifnone
       (A1 *> ZN) = (tphlh$A1$ZN,tplhl$A1$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OO01D2 (Z, A1, A2, B, C);
input  A1 ;
input  A2 ;
input  B ;
input  C ;
output Z ;

   or  (I0_out, A1, A2);
   and (I1_out, I0_out, B);
   or  (Z, I1_out, C);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$B$Z = 1.0,
       tphhl$B$Z = 1.0,
       tpllh$C$Z = 1.0,
       tphhl$C$Z = 1.0,
       tpllh$B$Z$A1_EQ_1_AN_A2_EQ_1_AN_C_EQ_0 = 1.0,
       tphhl$B$Z$A1_EQ_1_AN_A2_EQ_1_AN_C_EQ_0 = 1.0,
       tpllh$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_0 = 1.0,
       tphhl$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_0 = 1.0,
       tpllh$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_0 = 1.0,
       tphhl$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_0 = 1.0,
       tpllh$C$Z$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_0 = 1.0,
       tphhl$C$Z$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_0 = 1.0,
       tpllh$C$Z$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_0 = 1.0,
       tphhl$C$Z$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && B == 1'b0)
       (C *> Z) = (tpllh$C$Z$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_0, tphhl$C$Z$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b0)
       (C *> Z) = (tpllh$C$Z$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_0, tphhl$C$Z$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_0);
     ifnone
       (C *> Z) = (tpllh$C$Z,tphhl$C$Z);

     if (A1 == 1'b1 && A2 == 1'b1 && C == 1'b0)
       (B *> Z) = (tpllh$B$Z$A1_EQ_1_AN_A2_EQ_1_AN_C_EQ_0, tphhl$B$Z$A1_EQ_1_AN_A2_EQ_1_AN_C_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b0)
       (B *> Z) = (tpllh$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_0, tphhl$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b0)
       (B *> Z) = (tpllh$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_0, tphhl$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_0);
     ifnone
       (B *> Z) = (tpllh$B$Z,tphhl$B$Z);

     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OO01D4 (Z, A1, A2, B, C);
input  A1 ;
input  A2 ;
input  B ;
input  C ;
output Z ;

   or  (I0_out, A1, A2);
   and (I1_out, I0_out, B);
   or  (Z, I1_out, C);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$B$Z = 1.0,
       tphhl$B$Z = 1.0,
       tpllh$C$Z = 1.0,
       tphhl$C$Z = 1.0,
       tpllh$B$Z$A1_EQ_1_AN_A2_EQ_1_AN_C_EQ_0 = 1.0,
       tphhl$B$Z$A1_EQ_1_AN_A2_EQ_1_AN_C_EQ_0 = 1.0,
       tpllh$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_0 = 1.0,
       tphhl$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_0 = 1.0,
       tpllh$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_0 = 1.0,
       tphhl$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_0 = 1.0,
       tpllh$C$Z$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_0 = 1.0,
       tphhl$C$Z$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_0 = 1.0,
       tpllh$C$Z$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_0 = 1.0,
       tphhl$C$Z$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && B == 1'b0)
       (C *> Z) = (tpllh$C$Z$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_0, tphhl$C$Z$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b0)
       (C *> Z) = (tpllh$C$Z$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_0, tphhl$C$Z$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_0);
     ifnone
       (C *> Z) = (tpllh$C$Z,tphhl$C$Z);

     if (A1 == 1'b1 && A2 == 1'b1 && C == 1'b0)
       (B *> Z) = (tpllh$B$Z$A1_EQ_1_AN_A2_EQ_1_AN_C_EQ_0, tphhl$B$Z$A1_EQ_1_AN_A2_EQ_1_AN_C_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b0)
       (B *> Z) = (tpllh$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_0, tphhl$B$Z$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b0)
       (B *> Z) = (tpllh$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_0, tphhl$B$Z$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_0);
     ifnone
       (B *> Z) = (tpllh$B$Z,tphhl$B$Z);

     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OON1D1 (ZN, A1, A2, B, C);
input  A1 ;
input  A2 ;
input  B ;
input  C ;
output ZN ;

   or  (I0_out, A1, A2);
   and (I1_out, I0_out, B);
   or  (I2_out, I1_out, C);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$B$ZN = 1.0,
       tphlh$B$ZN = 1.0,
       tplhl$C$ZN = 1.0,
       tphlh$C$ZN = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_C_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_C_EQ_0 = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_0 = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_0 = 1.0,
       tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_0 = 1.0,
       tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_0 = 1.0,
       tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_0 = 1.0,
       tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && B == 1'b0)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_0, tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b0)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_0, tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_0);
     ifnone
       (C *> ZN) = (tphlh$C$ZN,tplhl$C$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && C == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_C_EQ_0, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_C_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_0, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_0, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_0);
     ifnone
       (B *> ZN) = (tphlh$B$ZN,tplhl$B$ZN);

     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OON1D2 (ZN, A1, A2, B, C);
input  A1 ;
input  A2 ;
input  B ;
input  C ;
output ZN ;

   or  (I0_out, A1, A2);
   and (I1_out, I0_out, B);
   or  (I2_out, I1_out, C);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$B$ZN = 1.0,
       tphlh$B$ZN = 1.0,
       tplhl$C$ZN = 1.0,
       tphlh$C$ZN = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_C_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_C_EQ_0 = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_0 = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_0 = 1.0,
       tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_0 = 1.0,
       tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_0 = 1.0,
       tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_0 = 1.0,
       tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && B == 1'b0)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_0, tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b0)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_0, tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_0);
     ifnone
       (C *> ZN) = (tphlh$C$ZN,tplhl$C$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && C == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_C_EQ_0, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_C_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_0, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_0, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_0);
     ifnone
       (B *> ZN) = (tphlh$B$ZN,tplhl$B$ZN);

     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OON1D4 (ZN, A1, A2, B, C);
input  A1 ;
input  A2 ;
input  B ;
input  C ;
output ZN ;

   or  (I0_out, A1, A2);
   and (I1_out, I0_out, B);
   or  (I2_out, I1_out, C);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tplhl$B$ZN = 1.0,
       tphlh$B$ZN = 1.0,
       tplhl$C$ZN = 1.0,
       tphlh$C$ZN = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_C_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_C_EQ_0 = 1.0,
       tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_0 = 1.0,
       tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_0 = 1.0,
       tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_0 = 1.0,
       tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_0 = 1.0,
       tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_0 = 1.0,
       tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_0 = 1.0,
       tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1 && B == 1'b0)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_0, tplhl$C$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b0)
       (C *> ZN) = (tphlh$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_0, tplhl$C$ZN$A1_EQ_0_AN_A2_EQ_0_AN_B_EQ_0);
     ifnone
       (C *> ZN) = (tphlh$C$ZN,tplhl$C$ZN);

     if (A1 == 1'b1 && A2 == 1'b1 && C == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_C_EQ_0, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_1_AN_C_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_0, tplhl$B$ZN$A1_EQ_1_AN_A2_EQ_0_AN_C_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b0)
       (B *> ZN) = (tphlh$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_0, tplhl$B$ZN$A1_EQ_0_AN_A2_EQ_1_AN_C_EQ_0);
     ifnone
       (B *> ZN) = (tphlh$B$ZN,tplhl$B$ZN);

     (A2 *> ZN) = (tphlh$A2$ZN, tplhl$A2$ZN);
     (A1 *> ZN) = (tphlh$A1$ZN, tplhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OR02D1 (Z, A1, A2);
input  A1 ;
input  A2 ;
output Z ;

   or  (Z, A1, A2);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0;

     // path delays
     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OR02D2 (Z, A1, A2);
input  A1 ;
input  A2 ;
output Z ;

   or  (Z, A1, A2);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0;

     // path delays
     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OR02D4 (Z, A1, A2);
input  A1 ;
input  A2 ;
output Z ;

   or  (Z, A1, A2);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0;

     // path delays
     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OR03D1 (Z, A1, A2, A3);
input  A1 ;
input  A2 ;
input  A3 ;
output Z ;

   or  (Z, A1, A2, A3);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$A3$Z = 1.0,
       tphhl$A3$Z = 1.0;

     // path delays
     (A3 *> Z) = (tpllh$A3$Z, tphhl$A3$Z);
     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OR03D2 (Z, A1, A2, A3);
input  A1 ;
input  A2 ;
input  A3 ;
output Z ;

   or  (Z, A1, A2, A3);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$A3$Z = 1.0,
       tphhl$A3$Z = 1.0;

     // path delays
     (A3 *> Z) = (tpllh$A3$Z, tphhl$A3$Z);
     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OR03D4 (Z, A1, A2, A3);
input  A1 ;
input  A2 ;
input  A3 ;
output Z ;

   or  (Z, A1, A2, A3);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$A3$Z = 1.0,
       tphhl$A3$Z = 1.0;

     // path delays
     (A3 *> Z) = (tpllh$A3$Z, tphhl$A3$Z);
     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OR04D1 (Z, A1, A2, A3, A4);
input  A1 ;
input  A2 ;
input  A3 ;
input  A4 ;
output Z ;

   or  (Z, A1, A2, A3, A4);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$A3$Z = 1.0,
       tphhl$A3$Z = 1.0,
       tpllh$A4$Z = 1.0,
       tphhl$A4$Z = 1.0;

     // path delays
     (A4 *> Z) = (tpllh$A4$Z, tphhl$A4$Z);
     (A3 *> Z) = (tpllh$A3$Z, tphhl$A3$Z);
     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OR04D2 (Z, A1, A2, A3, A4);
input  A1 ;
input  A2 ;
input  A3 ;
input  A4 ;
output Z ;

   or  (Z, A1, A2, A3, A4);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$A3$Z = 1.0,
       tphhl$A3$Z = 1.0,
       tpllh$A4$Z = 1.0,
       tphhl$A4$Z = 1.0;

     // path delays
     (A4 *> Z) = (tpllh$A4$Z, tphhl$A4$Z);
     (A3 *> Z) = (tpllh$A3$Z, tphhl$A3$Z);
     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OR04D4 (Z, A1, A2, A3, A4);
input  A1 ;
input  A2 ;
input  A3 ;
input  A4 ;
output Z ;

   or  (Z, A1, A2, A3, A4);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$A3$Z = 1.0,
       tphhl$A3$Z = 1.0,
       tpllh$A4$Z = 1.0,
       tphhl$A4$Z = 1.0;

     // path delays
     (A4 *> Z) = (tpllh$A4$Z, tphhl$A4$Z);
     (A3 *> Z) = (tpllh$A3$Z, tphhl$A3$Z);
     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OR06D2 (Z, A1, A2, A3, A4, A5, A6);
input  A1 ;
input  A2 ;
input  A3 ;
input  A4 ;
input  A5 ;
input  A6 ;
output Z ;

   or  (Z, A1, A2, A3, A4, A5, A6);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$A3$Z = 1.0,
       tphhl$A3$Z = 1.0,
       tpllh$A4$Z = 1.0,
       tphhl$A4$Z = 1.0,
       tpllh$A5$Z = 1.0,
       tphhl$A5$Z = 1.0,
       tpllh$A6$Z = 1.0,
       tphhl$A6$Z = 1.0;

     // path delays
     (A6 *> Z) = (tpllh$A6$Z, tphhl$A6$Z);
     (A5 *> Z) = (tpllh$A5$Z, tphhl$A5$Z);
     (A4 *> Z) = (tpllh$A4$Z, tphhl$A4$Z);
     (A3 *> Z) = (tpllh$A3$Z, tphhl$A3$Z);
     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OR06D4 (Z, A1, A2, A3, A4, A5, A6);
input  A1 ;
input  A2 ;
input  A3 ;
input  A4 ;
input  A5 ;
input  A6 ;
output Z ;

   or  (Z, A1, A2, A3, A4, A5, A6);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$A3$Z = 1.0,
       tphhl$A3$Z = 1.0,
       tpllh$A4$Z = 1.0,
       tphhl$A4$Z = 1.0,
       tpllh$A5$Z = 1.0,
       tphhl$A5$Z = 1.0,
       tpllh$A6$Z = 1.0,
       tphhl$A6$Z = 1.0;

     // path delays
     (A6 *> Z) = (tpllh$A6$Z, tphhl$A6$Z);
     (A5 *> Z) = (tpllh$A5$Z, tphhl$A5$Z);
     (A4 *> Z) = (tpllh$A4$Z, tphhl$A4$Z);
     (A3 *> Z) = (tpllh$A3$Z, tphhl$A3$Z);
     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OR08D2 (Z, A1, A2, A3, A4, A5, A6, A7, A8);
input  A1 ;
input  A2 ;
input  A3 ;
input  A4 ;
input  A5 ;
input  A6 ;
input  A7 ;
input  A8 ;
output Z ;

   or  (Z, A1, A2, A3, A4, A5, A6, A7, A8);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$A3$Z = 1.0,
       tphhl$A3$Z = 1.0,
       tpllh$A4$Z = 1.0,
       tphhl$A4$Z = 1.0,
       tpllh$A5$Z = 1.0,
       tphhl$A5$Z = 1.0,
       tpllh$A6$Z = 1.0,
       tphhl$A6$Z = 1.0,
       tpllh$A7$Z = 1.0,
       tphhl$A7$Z = 1.0,
       tpllh$A8$Z = 1.0,
       tphhl$A8$Z = 1.0;

     // path delays
     (A8 *> Z) = (tpllh$A8$Z, tphhl$A8$Z);
     (A7 *> Z) = (tpllh$A7$Z, tphhl$A7$Z);
     (A6 *> Z) = (tpllh$A6$Z, tphhl$A6$Z);
     (A5 *> Z) = (tpllh$A5$Z, tphhl$A5$Z);
     (A4 *> Z) = (tpllh$A4$Z, tphhl$A4$Z);
     (A3 *> Z) = (tpllh$A3$Z, tphhl$A3$Z);
     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OR08D4 (Z, A1, A2, A3, A4, A5, A6, A7, A8);
input  A1 ;
input  A2 ;
input  A3 ;
input  A4 ;
input  A5 ;
input  A6 ;
input  A7 ;
input  A8 ;
output Z ;

   or  (Z, A1, A2, A3, A4, A5, A6, A7, A8);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$A3$Z = 1.0,
       tphhl$A3$Z = 1.0,
       tpllh$A4$Z = 1.0,
       tphhl$A4$Z = 1.0,
       tpllh$A5$Z = 1.0,
       tphhl$A5$Z = 1.0,
       tpllh$A6$Z = 1.0,
       tphhl$A6$Z = 1.0,
       tpllh$A7$Z = 1.0,
       tphhl$A7$Z = 1.0,
       tpllh$A8$Z = 1.0,
       tphhl$A8$Z = 1.0;

     // path delays
     (A8 *> Z) = (tpllh$A8$Z, tphhl$A8$Z);
     (A7 *> Z) = (tpllh$A7$Z, tphhl$A7$Z);
     (A6 *> Z) = (tpllh$A6$Z, tphhl$A6$Z);
     (A5 *> Z) = (tpllh$A5$Z, tphhl$A5$Z);
     (A4 *> Z) = (tpllh$A4$Z, tphhl$A4$Z);
     (A3 *> Z) = (tpllh$A3$Z, tphhl$A3$Z);
     (A2 *> Z) = (tpllh$A2$Z, tphhl$A2$Z);
     (A1 *> Z) = (tpllh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OX01D1 (Z, A1, A2, B);
input  A1 ;
input  A2 ;
input  B ;
output Z ;

   or  (I0_out, A1, A2);
   xor (Z, I0_out, B);

   specify
     // delay parameters
    specparam
       tpllh$A1$Z = 1.0,
       tplhl$A1$Z = 1.0,
       tphlh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tplhl$A2$Z = 1.0,
       tphlh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$B$Z = 1.0,
       tplhl$B$Z = 1.0,
       tphlh$B$Z = 1.0,
       tphhl$B$Z = 1.0,
       tplhl$B$Z$A1_EQ_1_AN_A2_EQ_1 = 1.0,
       tphlh$B$Z$A1_EQ_1_AN_A2_EQ_1 = 1.0,
       tplhl$B$Z$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tphlh$B$Z$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tplhl$B$Z$A1_EQ_1_AN_A2_EQ_0 = 1.0,
       tphlh$B$Z$A1_EQ_1_AN_A2_EQ_0 = 1.0;

     // path delays
      (posedge B => (Z +: Z)) = (1.0, 1.0);
      (negedge B => (Z -: Z)) = (1.0, 1.0);

     if (A1 == 1'b1 && A2 == 1'b1)
       (B *> Z) = (tphlh$B$Z$A1_EQ_1_AN_A2_EQ_1, tplhl$B$Z$A1_EQ_1_AN_A2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0)
       (B *> Z) = (tphlh$B$Z$A1_EQ_1_AN_A2_EQ_0, tplhl$B$Z$A1_EQ_1_AN_A2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1)
       (B *> Z) = (tphlh$B$Z$A1_EQ_0_AN_A2_EQ_1, tplhl$B$Z$A1_EQ_0_AN_A2_EQ_1);
     /*   ifnone
       (B *> Z) = (tpllh$B$Z,tplhl$B$Z);

    (posedge B => (Z +: Z)) = (1.0, 1.0);
      (negedge B => (Z -: Z)) = (1.0, 1.0);
      if (A1 == 1'b1 && A2 == 1'b1) (B -=> Z) = (1.0, 1.0);
      if (A1 == 1'b0 && A2 == 1'b1) (B -=> Z) = (1.0, 1.0);
      if (A1 == 1'b1 && A2 == 1'b0) (B -=> Z) = (1.0, 1.0);*/
   

     (posedge A2 *> (Z +: !B)) = (tpllh$A2$Z, tplhl$A2$Z);
     (negedge A2 *> (Z +: B^A1)) = (tphlh$A2$Z, tphhl$A2$Z);
     (posedge A1 *> (Z +: !B)) = (tpllh$A1$Z, tplhl$A1$Z);
     (negedge A1 *> (Z +: B^A2)) = (tphlh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OX01D2 (Z, A1, A2, B);
input  A1 ;
input  A2 ;
input  B ;
output Z ;

   or  (I0_out, A1, A2);
   xor (Z, I0_out, B);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tplhl$A1$Z = 1.0,
       tphlh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tplhl$A2$Z = 1.0,
       tphlh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$B$Z = 1.0,
       tplhl$B$Z = 1.0,
       tphlh$B$Z = 1.0,
       tphhl$B$Z = 1.0,
       tplhl$B$Z$A1_EQ_1_AN_A2_EQ_1 = 1.0,
       tphlh$B$Z$A1_EQ_1_AN_A2_EQ_1 = 1.0,
       tplhl$B$Z$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tphlh$B$Z$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tplhl$B$Z$A1_EQ_1_AN_A2_EQ_0 = 1.0,
       tphlh$B$Z$A1_EQ_1_AN_A2_EQ_0 = 1.0;

     // path delays
      (posedge B => (Z +: Z)) = (1.0, 1.0);
      (negedge B => (Z -: Z)) = (1.0, 1.0);

     if (A1 == 1'b1 && A2 == 1'b1)
       (B *> Z) = (tphlh$B$Z$A1_EQ_1_AN_A2_EQ_1, tplhl$B$Z$A1_EQ_1_AN_A2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0)
       (B *> Z) = (tphlh$B$Z$A1_EQ_1_AN_A2_EQ_0, tplhl$B$Z$A1_EQ_1_AN_A2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1)
       (B *> Z) = (tphlh$B$Z$A1_EQ_0_AN_A2_EQ_1, tplhl$B$Z$A1_EQ_0_AN_A2_EQ_1);
 //    ifnone
   //    (B *> Z) = (tpllh$B$Z,tplhl$B$Z);

     (posedge A2 *> (Z +: !B)) = (tpllh$A2$Z, tplhl$A2$Z);
     (negedge A2 *> (Z +: B^A1)) = (tphlh$A2$Z, tphhl$A2$Z);
     (posedge A1 *> (Z +: !B)) = (tpllh$A1$Z, tplhl$A1$Z);
     (negedge A1 *> (Z +: B^A2)) = (tphlh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OX01D4 (Z, A1, A2, B);
input  A1 ;
input  A2 ;
input  B ;
output Z ;

   or  (I0_out, A1, A2);
   xor (Z, I0_out, B);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tplhl$A1$Z = 1.0,
       tphlh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tplhl$A2$Z = 1.0,
       tphlh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$B$Z = 1.0,
       tplhl$B$Z = 1.0,
       tphlh$B$Z = 1.0,
       tphhl$B$Z = 1.0,
       tplhl$B$Z$A1_EQ_1_AN_A2_EQ_1 = 1.0,
       tphlh$B$Z$A1_EQ_1_AN_A2_EQ_1 = 1.0,
       tplhl$B$Z$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tphlh$B$Z$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tplhl$B$Z$A1_EQ_1_AN_A2_EQ_0 = 1.0,
       tphlh$B$Z$A1_EQ_1_AN_A2_EQ_0 = 1.0;

     // path delays
      (posedge B => (Z +: Z)) = (1.0, 1.0);
      (negedge B => (Z -: Z)) = (1.0, 1.0);

     if (A1 == 1'b1 && A2 == 1'b1)
       (B *> Z) = (tphlh$B$Z$A1_EQ_1_AN_A2_EQ_1, tplhl$B$Z$A1_EQ_1_AN_A2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0)
       (B *> Z) = (tphlh$B$Z$A1_EQ_1_AN_A2_EQ_0, tplhl$B$Z$A1_EQ_1_AN_A2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1)
       (B *> Z) = (tphlh$B$Z$A1_EQ_0_AN_A2_EQ_1, tplhl$B$Z$A1_EQ_0_AN_A2_EQ_1);
 //    ifnone
   //    (B *> Z) = (tpllh$B$Z,tplhl$B$Z);

     (posedge A2 *> (Z +: !B)) = (tpllh$A2$Z, tplhl$A2$Z);
     (negedge A2 *> (Z +: B^A1)) = (tphlh$A2$Z, tphhl$A2$Z);
     (posedge A1 *> (Z +: !B)) = (tpllh$A1$Z, tplhl$A1$Z);
     (negedge A1 *> (Z +: B^A2)) = (tphlh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OX02D1 (Z, A1, A2, B1, B2);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
output Z ;

   or  (I0_out, A1, A2);
   or  (I1_out, B1, B2);
   xor (Z, I0_out, I1_out);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tplhl$A1$Z = 1.0,
       tphlh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tplhl$A2$Z = 1.0,
       tphlh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$B1$Z = 1.0,
       tplhl$B1$Z = 1.0,
       tphlh$B1$Z = 1.0,
       tphhl$B1$Z = 1.0,
       tpllh$B2$Z = 1.0,
       tplhl$B2$Z = 1.0,
       tphlh$B2$Z = 1.0,
       tphhl$B2$Z = 1.0,
       tplhl$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tphlh$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tplhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tphlh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tplhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0 = 1.0,
       tphlh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0 = 1.0;

     // path delays

      (posedge B2 => (Z +: Z)) = (1.0, 1.0);
      (negedge B2 => (Z -: Z)) = (1.0, 1.0);
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0)
       (B2 *> Z) = (tphlh$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0, tplhl$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
       (B2 *> Z) = (tphlh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0, tplhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
       (B2 *> Z) = (tphlh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0, tplhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0);
 //    ifnone
  //     (B2 *> Z) = (tpllh$B2$Z,tplhl$B2$Z);

      (posedge B1 => (Z +: Z)) = (1.0, 1.0);
      (negedge B1 => (Z -: Z)) = (1.0, 1.0);

     if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0)
       (B1 *> Z) = (tphlh$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0, tplhl$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
       (B1 *> Z) = (tphlh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0, tplhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
       (B1 *> Z) = (tphlh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0, tplhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0);
 //    ifnone
 //      (B1 *> Z) = (tpllh$B1$Z,tplhl$B1$Z);

      (posedge A2 => (Z +: Z)) = (1.0, 1.0);
      (negedge A2 => (Z -: Z)) = (1.0, 1.0);

     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (A2 *> Z) = (tphlh$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tplhl$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A2 *> Z) = (tphlh$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A2 *> Z) = (tphlh$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
  //   ifnone
  //     (A2 *> Z) = (tpllh$A2$Z,tplhl$A2$Z);

      (posedge A1 => (Z +: Z)) = (1.0, 1.0);
      (negedge A1 => (Z -: Z)) = (1.0, 1.0);

     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (A1 *> Z) = (tphlh$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tplhl$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A1 *> Z) = (tphlh$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A1 *> Z) = (tphlh$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
 //    ifnone
 //      (A1 *> Z) = (tpllh$A1$Z,tplhl$A1$Z);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OX02D2 (Z, A1, A2, B1, B2);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
output Z ;

   or  (I0_out, A1, A2);
   or  (I1_out, B1, B2);
   xor (Z, I0_out, I1_out);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tplhl$A1$Z = 1.0,
       tphlh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tplhl$A2$Z = 1.0,
       tphlh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$B1$Z = 1.0,
       tplhl$B1$Z = 1.0,
       tphlh$B1$Z = 1.0,
       tphhl$B1$Z = 1.0,
       tpllh$B2$Z = 1.0,
       tplhl$B2$Z = 1.0,
       tphlh$B2$Z = 1.0,
       tphhl$B2$Z = 1.0,
       tplhl$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tphlh$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tplhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tphlh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tplhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0 = 1.0,
       tphlh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0 = 1.0;

     // path delays
      (posedge B2 => (Z +: Z)) = (1.0, 1.0);
      (negedge B2 => (Z -: Z)) = (1.0, 1.0);
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0)
       (B2 *> Z) = (tphlh$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0, tplhl$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
       (B2 *> Z) = (tphlh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0, tplhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
       (B2 *> Z) = (tphlh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0, tplhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0);
  //   ifnone
   //    (B2 *> Z) = (tpllh$B2$Z,tplhl$B2$Z);

      (posedge B1 => (Z +: Z)) = (1.0, 1.0);
      (negedge B1 => (Z -: Z)) = (1.0, 1.0);

     if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0)
       (B1 *> Z) = (tphlh$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0, tplhl$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
       (B1 *> Z) = (tphlh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0, tplhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
       (B1 *> Z) = (tphlh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0, tplhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0);
//     ifnone
//       (B1 *> Z) = (tpllh$B1$Z,tplhl$B1$Z);

      (posedge A2 => (Z +: Z)) = (1.0, 1.0);
      (negedge A2 => (Z -: Z)) = (1.0, 1.0);

     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (A2 *> Z) = (tphlh$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tplhl$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A2 *> Z) = (tphlh$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A2 *> Z) = (tphlh$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
  //   ifnone
//       (A2 *> Z) = (tpllh$A2$Z,tplhl$A2$Z);

      (posedge A1 => (Z +: Z)) = (1.0, 1.0);
      (negedge A1 => (Z -: Z)) = (1.0, 1.0);

     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (A1 *> Z) = (tphlh$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tplhl$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A1 *> Z) = (tphlh$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A1 *> Z) = (tphlh$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
//     ifnone
//       (A1 *> Z) = (tpllh$A1$Z,tplhl$A1$Z);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OX02D4 (Z, A1, A2, B1, B2);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
output Z ;

   or  (I0_out, A1, A2);
   or  (I1_out, B1, B2);
   xor (Z, I0_out, I1_out);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tplhl$A1$Z = 1.0,
       tphlh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tplhl$A2$Z = 1.0,
       tphlh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$B1$Z = 1.0,
       tplhl$B1$Z = 1.0,
       tphlh$B1$Z = 1.0,
       tphhl$B1$Z = 1.0,
       tpllh$B2$Z = 1.0,
       tplhl$B2$Z = 1.0,
       tphlh$B2$Z = 1.0,
       tphhl$B2$Z = 1.0,
       tplhl$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphlh$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tplhl$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphlh$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tplhl$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tphlh$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tplhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0 = 1.0,
       tphlh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0 = 1.0,
       tplhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tphlh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tplhl$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tphlh$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tplhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0 = 1.0,
       tphlh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0 = 1.0;

     // path delays

      (posedge B2 => (Z +: Z)) = (1.0, 1.0);
      (negedge B2 => (Z -: Z)) = (1.0, 1.0);

     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0)
       (B2 *> Z) = (tphlh$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0, tplhl$B2$Z$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
       (B2 *> Z) = (tphlh$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0, tplhl$B2$Z$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
       (B2 *> Z) = (tphlh$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0, tplhl$B2$Z$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0);
    // ifnone
    //   (B2 *> Z) = (tpllh$B2$Z,tplhl$B2$Z);

      (posedge B1 => (Z +: Z)) = (1.0, 1.0);
      (negedge B1 => (Z -: Z)) = (1.0, 1.0);

     if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0)
       (B1 *> Z) = (tphlh$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0, tplhl$B1$Z$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
       (B1 *> Z) = (tphlh$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0, tplhl$B1$Z$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
       (B1 *> Z) = (tphlh$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0, tplhl$B1$Z$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0);
  //   ifnone
   //    (B1 *> Z) = (tpllh$B1$Z,tplhl$B1$Z);

      (posedge A2 => (Z +: Z)) = (1.0, 1.0);
      (negedge A2 => (Z -: Z)) = (1.0, 1.0);

     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (A2 *> Z) = (tphlh$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tplhl$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A2 *> Z) = (tphlh$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A2$Z$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A2 *> Z) = (tphlh$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A2$Z$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
  //   ifnone
  //     (A2 *> Z) = (tpllh$A2$Z,tplhl$A2$Z);

      (posedge A1 => (Z +: Z)) = (1.0, 1.0);
      (negedge A1 => (Z -: Z)) = (1.0, 1.0);

     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (A1 *> Z) = (tphlh$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tplhl$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A1 *> Z) = (tphlh$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tplhl$A1$Z$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A1 *> Z) = (tphlh$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tplhl$A1$Z$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
 //    ifnone
 //      (A1 *> Z) = (tpllh$A1$Z,tplhl$A1$Z);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OXN1D1 (ZN, A1, A2, B);
input  A1 ;
input  A2 ;
input  B ;
output ZN ;

   or  (I0_out, A1, A2);
   xor (I1_out, I0_out, B);
   not (ZN, I1_out);

   specify
     // delay parameters
     specparam
       tpllh$A1$ZN = 1.0,
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tphhl$A1$ZN = 1.0,
       tpllh$A2$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tphhl$A2$ZN = 1.0,
       tpllh$B$ZN = 1.0,
       tplhl$B$ZN = 1.0,
       tphlh$B$ZN = 1.0,
       tphhl$B$ZN = 1.0,
       tpllh$B$ZN$A1_EQ_1_AN_A2_EQ_1 = 1.0,
       tphhl$B$ZN$A1_EQ_1_AN_A2_EQ_1 = 1.0,
       tpllh$B$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tphhl$B$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tpllh$B$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0,
       tphhl$B$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0;

     // path delays
      (posedge B => (ZN +: ZN)) = (1.0, 1.0);
      (negedge B => (ZN -: ZN)) = (1.0, 1.0);


     if (A1 == 1'b1 && A2 == 1'b1)
       (B *> ZN) = (tpllh$B$ZN$A1_EQ_1_AN_A2_EQ_1, tphhl$B$ZN$A1_EQ_1_AN_A2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0)
       (B *> ZN) = (tpllh$B$ZN$A1_EQ_1_AN_A2_EQ_0, tphhl$B$ZN$A1_EQ_1_AN_A2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1)
       (B *> ZN) = (tpllh$B$ZN$A1_EQ_0_AN_A2_EQ_1, tphhl$B$ZN$A1_EQ_0_AN_A2_EQ_1);
//     ifnone
  //     (B *> ZN) = (tpllh$B$ZN,tplhl$B$ZN);

     (posedge A2 *> (ZN +: B)) = (tpllh$A2$ZN, tplhl$A2$ZN);
     (negedge A2 *> (ZN +: !(B^A1))) = (tphlh$A2$ZN, tphhl$A2$ZN);
     (posedge A1 *> (ZN +: B)) = (tpllh$A1$ZN, tplhl$A1$ZN);
     (negedge A1 *> (ZN +: !(B^A2))) = (tphlh$A1$ZN, tphhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OXN1D2 (ZN, A1, A2, B);
input  A1 ;
input  A2 ;
input  B ;
output ZN ;

   or  (I0_out, A1, A2);
   xor (I1_out, I0_out, B);
   not (ZN, I1_out);

   specify
     // delay parameters
     specparam
       tpllh$A1$ZN = 1.0,
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tphhl$A1$ZN = 1.0,
       tpllh$A2$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tphhl$A2$ZN = 1.0,
       tpllh$B$ZN = 1.0,
       tplhl$B$ZN = 1.0,
       tphlh$B$ZN = 1.0,
       tphhl$B$ZN = 1.0,
       tpllh$B$ZN$A1_EQ_1_AN_A2_EQ_1 = 1.0,
       tphhl$B$ZN$A1_EQ_1_AN_A2_EQ_1 = 1.0,
       tpllh$B$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tphhl$B$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tpllh$B$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0,
       tphhl$B$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0;

     // path delays

      (posedge B => (ZN +: ZN)) = (1.0, 1.0);
      (negedge B => (ZN -: ZN)) = (1.0, 1.0);

     if (A1 == 1'b1 && A2 == 1'b1)
       (B *> ZN) = (tpllh$B$ZN$A1_EQ_1_AN_A2_EQ_1, tphhl$B$ZN$A1_EQ_1_AN_A2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0)
       (B *> ZN) = (tpllh$B$ZN$A1_EQ_1_AN_A2_EQ_0, tphhl$B$ZN$A1_EQ_1_AN_A2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1)
       (B *> ZN) = (tpllh$B$ZN$A1_EQ_0_AN_A2_EQ_1, tphhl$B$ZN$A1_EQ_0_AN_A2_EQ_1);
 //    ifnone
   //    (B *> ZN) = (tpllh$B$ZN,tplhl$B$ZN);

     (posedge A2 *> (ZN +: B)) = (tpllh$A2$ZN, tplhl$A2$ZN);
     (negedge A2 *> (ZN +: !(B^A1))) = (tphlh$A2$ZN, tphhl$A2$ZN);
     (posedge A1 *> (ZN +: B)) = (tpllh$A1$ZN, tplhl$A1$ZN);
     (negedge A1 *> (ZN +: !(B^A2))) = (tphlh$A1$ZN, tphhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OXN1D4 (ZN, A1, A2, B);
input  A1 ;
input  A2 ;
input  B ;
output ZN ;

   or  (I0_out, A1, A2);
   xor (I1_out, I0_out, B);
   not (ZN, I1_out);

   specify
     // delay parameters
     specparam
       tpllh$A1$ZN = 1.0,
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tphhl$A1$ZN = 1.0,
       tpllh$A2$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tphhl$A2$ZN = 1.0,
       tpllh$B$ZN = 1.0,
       tplhl$B$ZN = 1.0,
       tphlh$B$ZN = 1.0,
       tphhl$B$ZN = 1.0,
       tpllh$B$ZN$A1_EQ_1_AN_A2_EQ_1 = 1.0,
       tphhl$B$ZN$A1_EQ_1_AN_A2_EQ_1 = 1.0,
       tpllh$B$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tphhl$B$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tpllh$B$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0,
       tphhl$B$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0;

     // path delays

      (posedge B => (ZN +: ZN)) = (1.0, 1.0);
      (negedge B => (ZN -: ZN)) = (1.0, 1.0);


     if (A1 == 1'b1 && A2 == 1'b1)
       (B *> ZN) = (tpllh$B$ZN$A1_EQ_1_AN_A2_EQ_1, tphhl$B$ZN$A1_EQ_1_AN_A2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0)
       (B *> ZN) = (tpllh$B$ZN$A1_EQ_1_AN_A2_EQ_0, tphhl$B$ZN$A1_EQ_1_AN_A2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1)
       (B *> ZN) = (tpllh$B$ZN$A1_EQ_0_AN_A2_EQ_1, tphhl$B$ZN$A1_EQ_0_AN_A2_EQ_1);
//     ifnone
  //     (B *> ZN) = (tpllh$B$ZN,tplhl$B$ZN);

     (posedge A2 *> (ZN +: B)) = (tpllh$A2$ZN, tplhl$A2$ZN);
     (negedge A2 *> (ZN +: !(B^A1))) = (tphlh$A2$ZN, tphhl$A2$ZN);
     (posedge A1 *> (ZN +: B)) = (tpllh$A1$ZN, tplhl$A1$ZN);
     (negedge A1 *> (ZN +: !(B^A2))) = (tphlh$A1$ZN, tphhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OXN2D1 (ZN, A1, A2, B1, B2);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
output ZN ;

   or  (I0_out, A1, A2);
   or  (I1_out, B1, B2);
   xor (I2_out, I0_out, I1_out);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tpllh$A1$ZN = 1.0,
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tphhl$A1$ZN = 1.0,
       tpllh$A2$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tphhl$A2$ZN = 1.0,
       tpllh$B1$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tphhl$B1$ZN = 1.0,
       tpllh$B2$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tphhl$B2$ZN = 1.0,
       tpllh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tpllh$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tpllh$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0 = 1.0,
       tpllh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0 = 1.0,
       tphhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0 = 1.0,
       tpllh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tphhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tpllh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tphhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0;

     // path delays
      (posedge B2 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge B2 => (ZN -: ZN)) = (1.0, 1.0);

     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0)
       (B2 *> ZN) = (tpllh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0, tphhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
       (B2 *> ZN) = (tpllh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0, tphhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
       (B2 *> ZN) = (tpllh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0, tphhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0);
 //    ifnone
 //      (B2 *> ZN) = (tpllh$B2$ZN,tplhl$B2$ZN);

      (posedge B1 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge B1 => (ZN -: ZN)) = (1.0, 1.0);

     if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0)
       (B1 *> ZN) = (tpllh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0, tphhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
       (B1 *> ZN) = (tpllh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0, tphhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
       (B1 *> ZN) = (tpllh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0, tphhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0);
  //   ifnone
  //     (B1 *> ZN) = (tpllh$B1$ZN,tplhl$B1$ZN);

      (posedge A2 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge A2 => (ZN -: ZN)) = (1.0, 1.0);

     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (A2 *> ZN) = (tpllh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tphhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A2 *> ZN) = (tpllh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A2 *> ZN) = (tpllh$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
  //   ifnone
  //     (A2 *> ZN) = (tpllh$A2$ZN,tplhl$A2$ZN);

      (posedge A1 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge A1 => (ZN -: ZN)) = (1.0, 1.0);

     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (A1 *> ZN) = (tpllh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tphhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A1 *> ZN) = (tpllh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A1 *> ZN) = (tpllh$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
   //  ifnone
   //    (A1 *> ZN) = (tpllh$A1$ZN,tplhl$A1$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OXN2D2 (ZN, A1, A2, B1, B2);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
output ZN ;

   or  (I0_out, A1, A2);
   or  (I1_out, B1, B2);
   xor (I2_out, I0_out, I1_out);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tpllh$A1$ZN = 1.0,
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tphhl$A1$ZN = 1.0,
       tpllh$A2$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tphhl$A2$ZN = 1.0,
       tpllh$B1$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tphhl$B1$ZN = 1.0,
       tpllh$B2$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tphhl$B2$ZN = 1.0,
       tpllh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tpllh$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tpllh$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0 = 1.0,
       tpllh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0 = 1.0,
       tphhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0 = 1.0,
       tpllh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tphhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tpllh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tphhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0;

     // path delays
      (posedge B2 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge B2 => (ZN -: ZN)) = (1.0, 1.0);

     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0)
       (B2 *> ZN) = (tpllh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0, tphhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
       (B2 *> ZN) = (tpllh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0, tphhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
       (B2 *> ZN) = (tpllh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0, tphhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0);
  //   ifnone
   //    (B2 *> ZN) = (tpllh$B2$ZN,tplhl$B2$ZN);

      (posedge B1 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge B1 => (ZN -: ZN)) = (1.0, 1.0);

     if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0)
       (B1 *> ZN) = (tpllh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0, tphhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
       (B1 *> ZN) = (tpllh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0, tphhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
       (B1 *> ZN) = (tpllh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0, tphhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0);
   //  ifnone
 //      (B1 *> ZN) = (tpllh$B1$ZN,tplhl$B1$ZN);

      (posedge A2 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge A2 => (ZN -: ZN)) = (1.0, 1.0);

     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (A2 *> ZN) = (tpllh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tphhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A2 *> ZN) = (tpllh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A2 *> ZN) = (tpllh$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
 //    ifnone
 //      (A2 *> ZN) = (tpllh$A2$ZN,tplhl$A2$ZN);

      (posedge A1 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge A1 => (ZN -: ZN)) = (1.0, 1.0);

     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (A1 *> ZN) = (tpllh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tphhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A1 *> ZN) = (tpllh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A1 *> ZN) = (tpllh$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
   //  ifnone
  //     (A1 *> ZN) = (tpllh$A1$ZN,tplhl$A1$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_OXN2D4 (ZN, A1, A2, B1, B2);
input  A1 ;
input  A2 ;
input  B1 ;
input  B2 ;
output ZN ;

   or  (I0_out, A1, A2);
   or  (I1_out, B1, B2);
   xor (I2_out, I0_out, I1_out);
   not (ZN, I2_out);

   specify
     // delay parameters
     specparam
       tpllh$A1$ZN = 1.0,
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tphhl$A1$ZN = 1.0,
       tpllh$A2$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tphhl$A2$ZN = 1.0,
       tpllh$B1$ZN = 1.0,
       tplhl$B1$ZN = 1.0,
       tphlh$B1$ZN = 1.0,
       tphhl$B1$ZN = 1.0,
       tpllh$B2$ZN = 1.0,
       tplhl$B2$ZN = 1.0,
       tphlh$B2$ZN = 1.0,
       tphhl$B2$ZN = 1.0,
       tpllh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tpllh$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tphhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1 = 1.0,
       tpllh$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tphhl$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1 = 1.0,
       tpllh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tphhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0 = 1.0,
       tpllh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0 = 1.0,
       tphhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0 = 1.0,
       tpllh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tphhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tpllh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tphhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0 = 1.0,
       tpllh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0 = 1.0,
       tphhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0 = 1.0;

     // path delays

      (posedge B2 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge B2 => (ZN -: ZN)) = (1.0, 1.0);
     if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0)
       (B2 *> ZN) = (tpllh$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0, tphhl$B2$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B1_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
       (B2 *> ZN) = (tpllh$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0, tphhl$B2$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B1_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
       (B2 *> ZN) = (tpllh$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0, tphhl$B2$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B1_EQ_0);
   //  ifnone
   //    (B2 *> ZN) = (tpllh$B2$ZN,tplhl$B2$ZN);

      (posedge B1 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge B1 => (ZN -: ZN)) = (1.0, 1.0);
     if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0)
       (B1 *> ZN) = (tpllh$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0, tphhl$B1$ZN$A1_EQ_1_AN_A2_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
       (B1 *> ZN) = (tpllh$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0, tphhl$B1$ZN$A1_EQ_1_AN_A2_EQ_0_AN_B2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
       (B1 *> ZN) = (tpllh$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0, tphhl$B1$ZN$A1_EQ_0_AN_A2_EQ_1_AN_B2_EQ_0);
  //   ifnone
  //     (B1 *> ZN) = (tpllh$B1$ZN,tplhl$B1$ZN);

      (posedge A2 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge A2 => (ZN -: ZN)) = (1.0, 1.0);
     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (A2 *> ZN) = (tpllh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tphhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A2 *> ZN) = (tpllh$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A2$ZN$A1_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A2 *> ZN) = (tpllh$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A2$ZN$A1_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
 //    ifnone
  //     (A2 *> ZN) = (tpllh$A2$ZN,tplhl$A2$ZN);

      (posedge A1 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge A1 => (ZN -: ZN)) = (1.0, 1.0);
     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
       (A1 *> ZN) = (tpllh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1, tphhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_1);
     if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
       (A1 *> ZN) = (tpllh$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0, tphhl$A1$ZN$A2_EQ_0_AN_B1_EQ_1_AN_B2_EQ_0);
     if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
       (A1 *> ZN) = (tpllh$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1, tphhl$A1$ZN$A2_EQ_0_AN_B1_EQ_0_AN_B2_EQ_1);
 //    ifnone
 //      (A1 *> ZN) = (tpllh$A1$ZN,tplhl$A1$ZN);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_SDF01D1 (Q, QN, CP, D, SE, SI);
input  CP ;
input  D ;
input  SE ;
input  SI ;
output Q ;
output QN ;
reg NOTIFIER ;
reg ReSeT;

`ifdef  RSTn_lib
	 initial begin
		ReSeT = 0 ;
		#3 ReSeT = 1 ;
		#111 ReSeT = 0 ;
	end
  `else initial  ReSeT = 0;
`endif


   udp_dff (N_S_XM27_G, I0_D, CP, ReSeT , 1'B0, NOTIFIER);


   udp_mux2 (I0_D, D, SI, SE);
   not (N_NET0130_XM24_D, N_S_XM27_G);
   buf (Q, N_S_XM27_G);
   not (QN, N_S_XM27_G);
   not (I7_out, D);
   and (D_EQ_0_AN_SI_EQ_1, I7_out, SI);
   not (I9_out, SI);
   and (D_EQ_1_AN_SI_EQ_0, D, I9_out);
   not (I11_out, D);
   not (I12_out, SE);
   not (I14_out, SI);
   and (D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, I11_out, I12_out, I14_out);

   specify
     // delay parameters
     specparam
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tpllh$CP$QN = 1.0,
       tplhl$CP$QN = 1.0,
       tminpwh$CP$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwl$CP$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tsetup_negedge$D$CP$SE_EQ_0 = 1.0,
       thold_negedge$D$CP$SE_EQ_0 = 1.0,
       tsetup_negedge$SE$CP$D_EQ_0_AN_SI_EQ_1 = 1.0,
       thold_negedge$SE$CP$D_EQ_0_AN_SI_EQ_1 = 1.0,
       tsetup_negedge$SE$CP$D_EQ_1_AN_SI_EQ_0 = 1.0,
       thold_negedge$SE$CP$D_EQ_1_AN_SI_EQ_0 = 1.0,
       tsetup_negedge$SI$CP$SE_EQ_1 = 1.0,
       thold_negedge$SI$CP$SE_EQ_1 = 1.0,
       tsetup_posedge$D$CP$SE_EQ_0 = 1.0,
       thold_posedge$D$CP$SE_EQ_0 = 1.0,
       tsetup_posedge$SE$CP$D_EQ_0_AN_SI_EQ_1 = 1.0,
       thold_posedge$SE$CP$D_EQ_0_AN_SI_EQ_1 = 1.0,
       tsetup_posedge$SE$CP$D_EQ_1_AN_SI_EQ_0 = 1.0,
       thold_posedge$SE$CP$D_EQ_1_AN_SI_EQ_0 = 1.0,
       tsetup_posedge$SI$CP$SE_EQ_1 = 1.0,
       thold_posedge$SI$CP$SE_EQ_1 = 1.0;

     // path delays
     (posedge CP *> (QN -: SE?SI:D)) = (tpllh$CP$QN, tplhl$CP$QN);
     (posedge CP *> (Q +: SE?SI:D)) = (tpllh$CP$Q, tplhl$CP$Q);
     $setuphold(posedge CP &&& SE == 1'b0, negedge D, tsetup_negedge$D$CP$SE_EQ_0, thold_negedge$D$CP$SE_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& D_EQ_0_AN_SI_EQ_1 == 1'b1, negedge SE, tsetup_negedge$SE$CP$D_EQ_0_AN_SI_EQ_1, thold_negedge$SE$CP$D_EQ_0_AN_SI_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& D_EQ_1_AN_SI_EQ_0 == 1'b1, negedge SE, tsetup_negedge$SE$CP$D_EQ_1_AN_SI_EQ_0, thold_negedge$SE$CP$D_EQ_1_AN_SI_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& SE == 1'b1, negedge SI, tsetup_negedge$SI$CP$SE_EQ_1, thold_negedge$SI$CP$SE_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& SE == 1'b0, posedge D, tsetup_posedge$D$CP$SE_EQ_0, thold_posedge$D$CP$SE_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& D_EQ_0_AN_SI_EQ_1 == 1'b1, posedge SE, tsetup_posedge$SE$CP$D_EQ_0_AN_SI_EQ_1, thold_posedge$SE$CP$D_EQ_0_AN_SI_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& D_EQ_1_AN_SI_EQ_0 == 1'b1, posedge SE, tsetup_posedge$SE$CP$D_EQ_1_AN_SI_EQ_0, thold_posedge$SE$CP$D_EQ_1_AN_SI_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& SE == 1'b1, posedge SI, tsetup_posedge$SI$CP$SE_EQ_1, thold_posedge$SI$CP$SE_EQ_1, NOTIFIER);
     $width(posedge CP &&& D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwh$CP$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(negedge CP &&& D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$CP$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_SDF01D2 (Q, QN, CP, D, SE, SI);
input  CP ;
input  D ;
input  SE ;
input  SI ;
output Q ;
output QN ;
reg NOTIFIER ;
reg ReSeT;

`ifdef  RSTn_lib
	 initial begin
		ReSeT = 0 ;
		#3 ReSeT = 1 ;
		#111 ReSeT = 0 ;
	end
  `else initial  ReSeT = 0;
`endif

   udp_mux2 (I0_D, D, SI, SE);
   udp_dff (N_S_XM27_G, I0_D, CP, ReSeT , 1'B0, NOTIFIER);
   not (N_NET0130_XM24_D, N_S_XM27_G);
   buf (Q, N_S_XM27_G);
   not (QN, N_S_XM27_G);
   not (I7_out, D);
   and (D_EQ_0_AN_SI_EQ_1, I7_out, SI);
   not (I9_out, SI);
   and (D_EQ_1_AN_SI_EQ_0, D, I9_out);
   not (I11_out, D);
   not (I12_out, SE);
   not (I14_out, SI);
   and (D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, I11_out, I12_out, I14_out);

   specify
     // delay parameters
     specparam
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tpllh$CP$QN = 1.0,
       tplhl$CP$QN = 1.0,
       tminpwh$CP$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwl$CP$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tsetup_negedge$D$CP$SE_EQ_0 = 1.0,
       thold_negedge$D$CP$SE_EQ_0 = 1.0,
       tsetup_negedge$SE$CP$D_EQ_0_AN_SI_EQ_1 = 1.0,
       thold_negedge$SE$CP$D_EQ_0_AN_SI_EQ_1 = 1.0,
       tsetup_negedge$SE$CP$D_EQ_1_AN_SI_EQ_0 = 1.0,
       thold_negedge$SE$CP$D_EQ_1_AN_SI_EQ_0 = 1.0,
       tsetup_negedge$SI$CP$SE_EQ_1 = 1.0,
       thold_negedge$SI$CP$SE_EQ_1 = 1.0,
       tsetup_posedge$D$CP$SE_EQ_0 = 1.0,
       thold_posedge$D$CP$SE_EQ_0 = 1.0,
       tsetup_posedge$SE$CP$D_EQ_0_AN_SI_EQ_1 = 1.0,
       thold_posedge$SE$CP$D_EQ_0_AN_SI_EQ_1 = 1.0,
       tsetup_posedge$SE$CP$D_EQ_1_AN_SI_EQ_0 = 1.0,
       thold_posedge$SE$CP$D_EQ_1_AN_SI_EQ_0 = 1.0,
       tsetup_posedge$SI$CP$SE_EQ_1 = 1.0,
       thold_posedge$SI$CP$SE_EQ_1 = 1.0;

     // path delays
     (posedge CP *> (QN -: SE?SI:D)) = (tpllh$CP$QN, tplhl$CP$QN);
     (posedge CP *> (Q +: SE?SI:D)) = (tpllh$CP$Q, tplhl$CP$Q);
     $setuphold(posedge CP &&& SE == 1'b0, negedge D, tsetup_negedge$D$CP$SE_EQ_0, thold_negedge$D$CP$SE_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& D_EQ_0_AN_SI_EQ_1 == 1'b1, negedge SE, tsetup_negedge$SE$CP$D_EQ_0_AN_SI_EQ_1, thold_negedge$SE$CP$D_EQ_0_AN_SI_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& D_EQ_1_AN_SI_EQ_0 == 1'b1, negedge SE, tsetup_negedge$SE$CP$D_EQ_1_AN_SI_EQ_0, thold_negedge$SE$CP$D_EQ_1_AN_SI_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& SE == 1'b1, negedge SI, tsetup_negedge$SI$CP$SE_EQ_1, thold_negedge$SI$CP$SE_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& SE == 1'b0, posedge D, tsetup_posedge$D$CP$SE_EQ_0, thold_posedge$D$CP$SE_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& D_EQ_0_AN_SI_EQ_1 == 1'b1, posedge SE, tsetup_posedge$SE$CP$D_EQ_0_AN_SI_EQ_1, thold_posedge$SE$CP$D_EQ_0_AN_SI_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& D_EQ_1_AN_SI_EQ_0 == 1'b1, posedge SE, tsetup_posedge$SE$CP$D_EQ_1_AN_SI_EQ_0, thold_posedge$SE$CP$D_EQ_1_AN_SI_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& SE == 1'b1, posedge SI, tsetup_posedge$SI$CP$SE_EQ_1, thold_posedge$SI$CP$SE_EQ_1, NOTIFIER);
     $width(posedge CP &&& D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwh$CP$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(negedge CP &&& D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$CP$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_SDF01D4 (Q, QN, CP, D, SE, SI);
input  CP ;
input  D ;
input  SE ;
input  SI ;
output Q ;
output QN ;
reg NOTIFIER ;
reg ReSeT;

`ifdef  RSTn_lib
	 initial begin
		ReSeT = 0 ;
		#3 ReSeT = 1 ;
		#111 ReSeT = 0 ;
	end
  `else initial  ReSeT = 0;
`endif


   udp_mux2 (I0_D, D, SI, SE);
   udp_dff (N_S_XM27_G, I0_D, CP, ReSeT, 1'B0, NOTIFIER);
   not (N_NET0130_XM24_D, N_S_XM27_G);
   buf (Q, N_S_XM27_G);
   not (QN, N_S_XM27_G);
   not (I7_out, D);
   and (D_EQ_0_AN_SI_EQ_1, I7_out, SI);
   not (I9_out, SI);
   and (D_EQ_1_AN_SI_EQ_0, D, I9_out);
   not (I11_out, D);
   not (I12_out, SE);
   not (I14_out, SI);
   and (D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, I11_out, I12_out, I14_out);

   specify
     // delay parameters
     specparam
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tpllh$CP$QN = 1.0,
       tplhl$CP$QN = 1.0,
       tminpwh$CP$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwl$CP$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tsetup_negedge$D$CP$SE_EQ_0 = 1.0,
       thold_negedge$D$CP$SE_EQ_0 = 1.0,
       tsetup_negedge$SE$CP$D_EQ_0_AN_SI_EQ_1 = 1.0,
       thold_negedge$SE$CP$D_EQ_0_AN_SI_EQ_1 = 1.0,
       tsetup_negedge$SE$CP$D_EQ_1_AN_SI_EQ_0 = 1.0,
       thold_negedge$SE$CP$D_EQ_1_AN_SI_EQ_0 = 1.0,
       tsetup_negedge$SI$CP$SE_EQ_1 = 1.0,
       thold_negedge$SI$CP$SE_EQ_1 = 1.0,
       tsetup_posedge$D$CP$SE_EQ_0 = 1.0,
       thold_posedge$D$CP$SE_EQ_0 = 1.0,
       tsetup_posedge$SE$CP$D_EQ_0_AN_SI_EQ_1 = 1.0,
       thold_posedge$SE$CP$D_EQ_0_AN_SI_EQ_1 = 1.0,
       tsetup_posedge$SE$CP$D_EQ_1_AN_SI_EQ_0 = 1.0,
       thold_posedge$SE$CP$D_EQ_1_AN_SI_EQ_0 = 1.0,
       tsetup_posedge$SI$CP$SE_EQ_1 = 1.0,
       thold_posedge$SI$CP$SE_EQ_1 = 1.0;

     // path delays
     (posedge CP *> (QN -: SE?SI:D)) = (tpllh$CP$QN, tplhl$CP$QN);
     (posedge CP *> (Q +: SE?SI:D)) = (tpllh$CP$Q, tplhl$CP$Q);
     $setuphold(posedge CP &&& SE == 1'b0, negedge D, tsetup_negedge$D$CP$SE_EQ_0, thold_negedge$D$CP$SE_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& D_EQ_0_AN_SI_EQ_1 == 1'b1, negedge SE, tsetup_negedge$SE$CP$D_EQ_0_AN_SI_EQ_1, thold_negedge$SE$CP$D_EQ_0_AN_SI_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& D_EQ_1_AN_SI_EQ_0 == 1'b1, negedge SE, tsetup_negedge$SE$CP$D_EQ_1_AN_SI_EQ_0, thold_negedge$SE$CP$D_EQ_1_AN_SI_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& SE == 1'b1, negedge SI, tsetup_negedge$SI$CP$SE_EQ_1, thold_negedge$SI$CP$SE_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& SE == 1'b0, posedge D, tsetup_posedge$D$CP$SE_EQ_0, thold_posedge$D$CP$SE_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& D_EQ_0_AN_SI_EQ_1 == 1'b1, posedge SE, tsetup_posedge$SE$CP$D_EQ_0_AN_SI_EQ_1, thold_posedge$SE$CP$D_EQ_0_AN_SI_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& D_EQ_1_AN_SI_EQ_0 == 1'b1, posedge SE, tsetup_posedge$SE$CP$D_EQ_1_AN_SI_EQ_0, thold_posedge$SE$CP$D_EQ_1_AN_SI_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& SE == 1'b1, posedge SI, tsetup_posedge$SI$CP$SE_EQ_1, thold_posedge$SI$CP$SE_EQ_1, NOTIFIER);
     $width(posedge CP &&& D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwh$CP$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(negedge CP &&& D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$CP$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_SDF02D1 (Q, QN, CDN, CP, D, SE, SI);
input  CDN ;
input  CP ;
input  D ;
input  SE ;
input  SI ;
output Q ;
output QN ;
reg NOTIFIER ;

   udp_mux2 (I0_D, D, SI, SE);
   not (I0_CLEAR, CDN);
   udp_dff (N_S_XM31_G, I0_D, CP, I0_CLEAR, 1'B0, NOTIFIER);
   not (N_NET0130_XM28_D, N_S_XM31_G);
   buf (Q, N_S_XM31_G);
   not (QN, N_S_XM31_G);
   and (CDN_EQ_1_AN_SE_EQ_1, CDN, SE);
   not (I9_out, SE);
   and (CDN_EQ_1_AN_SE_EQ_0, CDN, I9_out);
   not (I11_out, D);
   and (D_EQ_0_AN_SE_EQ_1_AN_SI_EQ_1, I11_out, SE, SI);
   not (I14_out, D);
   not (I15_out, SE);
   not (I17_out, SI);
   and (D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, I14_out, I15_out, I17_out);
   not (I19_out, D);
   not (I21_out, SE);
   not (I23_out, SI);
   and (CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, CDN, I19_out, I21_out, I23_out);

   specify
     // delay parameters
     specparam
       tphhl$CDN$Q = 1.0,
       tphlh$CDN$QN = 1.0,
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tpllh$CP$QN = 1.0,
       tplhl$CP$QN = 1.0,
       tminpwl$CDN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwh$CP$CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwl$CP$CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tsetup_negedge$D$CP$CDN_EQ_1_AN_SE_EQ_0 = 1.0,
       thold_negedge$D$CP$CDN_EQ_1_AN_SE_EQ_0 = 1.0,
       tsetup_negedge$SE$CP$CDN_EQ_1 = 1.0,
       thold_negedge$SE$CP$CDN_EQ_1 = 1.0,
       tsetup_negedge$SI$CP$CDN_EQ_1_AN_SE_EQ_1 = 1.0,
       thold_negedge$SI$CP$CDN_EQ_1_AN_SE_EQ_1 = 1.0,
       tsetup_posedge$D$CP$CDN_EQ_1_AN_SE_EQ_0 = 1.0,
       thold_posedge$D$CP$CDN_EQ_1_AN_SE_EQ_0 = 1.0,
       tsetup_posedge$SE$CP$CDN_EQ_1 = 1.0,
       thold_posedge$SE$CP$CDN_EQ_1 = 1.0,
       tsetup_posedge$SI$CP$CDN_EQ_1_AN_SE_EQ_1 = 1.0,
       thold_posedge$SI$CP$CDN_EQ_1_AN_SE_EQ_1 = 1.0,
       trec$CDN$CP$D_EQ_0_AN_SE_EQ_1_AN_SI_EQ_1 = 1.0,
       trem$CDN$CP$D_EQ_0_AN_SE_EQ_1_AN_SI_EQ_1 = 1.0;

     // path delays
     (posedge CP *> (QN -: SE?SI:D)) = (tpllh$CP$QN, tplhl$CP$QN);
     (posedge CP *> (Q +: SE?SI:D)) = (tpllh$CP$Q, tplhl$CP$Q);
     (negedge CDN *> (QN +: 1'b1)) = (tphlh$CDN$QN, 0);
     (negedge CDN *> (Q -: 1'b1)) = (0, tphhl$CDN$Q);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_SE_EQ_0 == 1'b1, negedge D, tsetup_negedge$D$CP$CDN_EQ_1_AN_SE_EQ_0, thold_negedge$D$CP$CDN_EQ_1_AN_SE_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& CDN == 1'b1, negedge SE, tsetup_negedge$SE$CP$CDN_EQ_1, thold_negedge$SE$CP$CDN_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_SE_EQ_1 == 1'b1, negedge SI, tsetup_negedge$SI$CP$CDN_EQ_1_AN_SE_EQ_1, thold_negedge$SI$CP$CDN_EQ_1_AN_SE_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_SE_EQ_0 == 1'b1, posedge D, tsetup_posedge$D$CP$CDN_EQ_1_AN_SE_EQ_0, thold_posedge$D$CP$CDN_EQ_1_AN_SE_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& CDN == 1'b1, posedge SE, tsetup_posedge$SE$CP$CDN_EQ_1, thold_posedge$SE$CP$CDN_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_SE_EQ_1 == 1'b1, posedge SI, tsetup_posedge$SI$CP$CDN_EQ_1_AN_SE_EQ_1, thold_posedge$SI$CP$CDN_EQ_1_AN_SE_EQ_1, NOTIFIER);
     $recrem(posedge CDN, posedge CP &&& D_EQ_0_AN_SE_EQ_1_AN_SI_EQ_1 == 1'b1, trec$CDN$CP$D_EQ_0_AN_SE_EQ_1_AN_SI_EQ_1, trem$CDN$CP$D_EQ_0_AN_SE_EQ_1_AN_SI_EQ_1, NOTIFIER);
     $width(negedge CDN &&& D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$CDN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(posedge CP &&& CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwh$CP$CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(negedge CP &&& CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$CP$CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_SDF02D2 (Q, QN, CDN, CP, D, SE, SI);
input  CDN ;
input  CP ;
input  D ;
input  SE ;
input  SI ;
output Q ;
output QN ;
reg NOTIFIER ;

   udp_mux2 (I0_D, D, SI, SE);
   not (I0_CLEAR, CDN);
   udp_dff (N_S_XM31_G, I0_D, CP, I0_CLEAR, 1'B0, NOTIFIER);
   not (N_NET0130_XM28_D, N_S_XM31_G);
   buf (Q, N_S_XM31_G);
   not (QN, N_S_XM31_G);
   and (CDN_EQ_1_AN_SE_EQ_1, CDN, SE);
   not (I9_out, SE);
   and (CDN_EQ_1_AN_SE_EQ_0, CDN, I9_out);
   not (I11_out, D);
   and (D_EQ_0_AN_SE_EQ_1_AN_SI_EQ_1, I11_out, SE, SI);
   not (I14_out, D);
   not (I15_out, SE);
   not (I17_out, SI);
   and (D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, I14_out, I15_out, I17_out);
   not (I19_out, D);
   not (I21_out, SE);
   not (I23_out, SI);
   and (CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, CDN, I19_out, I21_out, I23_out);

   specify
     // delay parameters
     specparam
       tphhl$CDN$Q = 1.0,
       tphlh$CDN$QN = 1.0,
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tpllh$CP$QN = 1.0,
       tplhl$CP$QN = 1.0,
       tminpwl$CDN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwh$CP$CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwl$CP$CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tsetup_negedge$D$CP$CDN_EQ_1_AN_SE_EQ_0 = 1.0,
       thold_negedge$D$CP$CDN_EQ_1_AN_SE_EQ_0 = 1.0,
       tsetup_negedge$SE$CP$CDN_EQ_1 = 1.0,
       thold_negedge$SE$CP$CDN_EQ_1 = 1.0,
       tsetup_negedge$SI$CP$CDN_EQ_1_AN_SE_EQ_1 = 1.0,
       thold_negedge$SI$CP$CDN_EQ_1_AN_SE_EQ_1 = 1.0,
       tsetup_posedge$D$CP$CDN_EQ_1_AN_SE_EQ_0 = 1.0,
       thold_posedge$D$CP$CDN_EQ_1_AN_SE_EQ_0 = 1.0,
       tsetup_posedge$SE$CP$CDN_EQ_1 = 1.0,
       thold_posedge$SE$CP$CDN_EQ_1 = 1.0,
       tsetup_posedge$SI$CP$CDN_EQ_1_AN_SE_EQ_1 = 1.0,
       thold_posedge$SI$CP$CDN_EQ_1_AN_SE_EQ_1 = 1.0,
       trec$CDN$CP$D_EQ_0_AN_SE_EQ_1_AN_SI_EQ_1 = 1.0,
       trem$CDN$CP$D_EQ_0_AN_SE_EQ_1_AN_SI_EQ_1 = 1.0;

     // path delays
     (posedge CP *> (QN -: SE?SI:D)) = (tpllh$CP$QN, tplhl$CP$QN);
     (posedge CP *> (Q +: SE?SI:D)) = (tpllh$CP$Q, tplhl$CP$Q);
     (negedge CDN *> (QN +: 1'b1)) = (tphlh$CDN$QN, 0);
     (negedge CDN *> (Q -: 1'b1)) = (0, tphhl$CDN$Q);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_SE_EQ_0 == 1'b1, negedge D, tsetup_negedge$D$CP$CDN_EQ_1_AN_SE_EQ_0, thold_negedge$D$CP$CDN_EQ_1_AN_SE_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& CDN == 1'b1, negedge SE, tsetup_negedge$SE$CP$CDN_EQ_1, thold_negedge$SE$CP$CDN_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_SE_EQ_1 == 1'b1, negedge SI, tsetup_negedge$SI$CP$CDN_EQ_1_AN_SE_EQ_1, thold_negedge$SI$CP$CDN_EQ_1_AN_SE_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_SE_EQ_0 == 1'b1, posedge D, tsetup_posedge$D$CP$CDN_EQ_1_AN_SE_EQ_0, thold_posedge$D$CP$CDN_EQ_1_AN_SE_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& CDN == 1'b1, posedge SE, tsetup_posedge$SE$CP$CDN_EQ_1, thold_posedge$SE$CP$CDN_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_SE_EQ_1 == 1'b1, posedge SI, tsetup_posedge$SI$CP$CDN_EQ_1_AN_SE_EQ_1, thold_posedge$SI$CP$CDN_EQ_1_AN_SE_EQ_1, NOTIFIER);
     $recrem(posedge CDN, posedge CP &&& D_EQ_0_AN_SE_EQ_1_AN_SI_EQ_1 == 1'b1, trec$CDN$CP$D_EQ_0_AN_SE_EQ_1_AN_SI_EQ_1, trem$CDN$CP$D_EQ_0_AN_SE_EQ_1_AN_SI_EQ_1, NOTIFIER);
     $width(negedge CDN &&& D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$CDN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(posedge CP &&& CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwh$CP$CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(negedge CP &&& CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$CP$CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_SDF02D4 (Q, QN, CDN, CP, D, SE, SI);
input  CDN ;
input  CP ;
input  D ;
input  SE ;
input  SI ;
output Q ;
output QN ;
reg NOTIFIER ;

   udp_mux2 (I0_D, D, SI, SE);
   not (I0_CLEAR, CDN);
   udp_dff (N_S_XM31_G, I0_D, CP, I0_CLEAR, 1'B0, NOTIFIER);
   not (N_NET0130_XM28_D, N_S_XM31_G);
   buf (Q, N_S_XM31_G);
   not (QN, N_S_XM31_G);
   and (CDN_EQ_1_AN_SE_EQ_1, CDN, SE);
   not (I9_out, SE);
   and (CDN_EQ_1_AN_SE_EQ_0, CDN, I9_out);
   not (I11_out, D);
   and (D_EQ_0_AN_SE_EQ_1_AN_SI_EQ_1, I11_out, SE, SI);
   not (I14_out, D);
   not (I15_out, SE);
   not (I17_out, SI);
   and (D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, I14_out, I15_out, I17_out);
   not (I19_out, D);
   not (I21_out, SE);
   not (I23_out, SI);
   and (CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, CDN, I19_out, I21_out, I23_out);

   specify
     // delay parameters
     specparam
       tphhl$CDN$Q = 1.0,
       tphlh$CDN$QN = 1.0,
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tpllh$CP$QN = 1.0,
       tplhl$CP$QN = 1.0,
       tminpwl$CDN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwh$CP$CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwl$CP$CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tsetup_negedge$D$CP$CDN_EQ_1_AN_SE_EQ_0 = 1.0,
       thold_negedge$D$CP$CDN_EQ_1_AN_SE_EQ_0 = 1.0,
       tsetup_negedge$SE$CP$CDN_EQ_1 = 1.0,
       thold_negedge$SE$CP$CDN_EQ_1 = 1.0,
       tsetup_negedge$SI$CP$CDN_EQ_1_AN_SE_EQ_1 = 1.0,
       thold_negedge$SI$CP$CDN_EQ_1_AN_SE_EQ_1 = 1.0,
       tsetup_posedge$D$CP$CDN_EQ_1_AN_SE_EQ_0 = 1.0,
       thold_posedge$D$CP$CDN_EQ_1_AN_SE_EQ_0 = 1.0,
       tsetup_posedge$SE$CP$CDN_EQ_1 = 1.0,
       thold_posedge$SE$CP$CDN_EQ_1 = 1.0,
       tsetup_posedge$SI$CP$CDN_EQ_1_AN_SE_EQ_1 = 1.0,
       thold_posedge$SI$CP$CDN_EQ_1_AN_SE_EQ_1 = 1.0,
       trec$CDN$CP$D_EQ_0_AN_SE_EQ_1_AN_SI_EQ_1 = 1.0,
       trem$CDN$CP$D_EQ_0_AN_SE_EQ_1_AN_SI_EQ_1 = 1.0;

     // path delays
     (posedge CP *> (QN -: SE?SI:D)) = (tpllh$CP$QN, tplhl$CP$QN);
     (posedge CP *> (Q +: SE?SI:D)) = (tpllh$CP$Q, tplhl$CP$Q);
     (negedge CDN *> (QN +: 1'b1)) = (tphlh$CDN$QN, 0);
     (negedge CDN *> (Q -: 1'b1)) = (0, tphhl$CDN$Q);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_SE_EQ_0 == 1'b1, negedge D, tsetup_negedge$D$CP$CDN_EQ_1_AN_SE_EQ_0, thold_negedge$D$CP$CDN_EQ_1_AN_SE_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& CDN == 1'b1, negedge SE, tsetup_negedge$SE$CP$CDN_EQ_1, thold_negedge$SE$CP$CDN_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_SE_EQ_1 == 1'b1, negedge SI, tsetup_negedge$SI$CP$CDN_EQ_1_AN_SE_EQ_1, thold_negedge$SI$CP$CDN_EQ_1_AN_SE_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_SE_EQ_0 == 1'b1, posedge D, tsetup_posedge$D$CP$CDN_EQ_1_AN_SE_EQ_0, thold_posedge$D$CP$CDN_EQ_1_AN_SE_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& CDN == 1'b1, posedge SE, tsetup_posedge$SE$CP$CDN_EQ_1, thold_posedge$SE$CP$CDN_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_SE_EQ_1 == 1'b1, posedge SI, tsetup_posedge$SI$CP$CDN_EQ_1_AN_SE_EQ_1, thold_posedge$SI$CP$CDN_EQ_1_AN_SE_EQ_1, NOTIFIER);
     $recrem(posedge CDN, posedge CP &&& D_EQ_0_AN_SE_EQ_1_AN_SI_EQ_1 == 1'b1, trec$CDN$CP$D_EQ_0_AN_SE_EQ_1_AN_SI_EQ_1, trem$CDN$CP$D_EQ_0_AN_SE_EQ_1_AN_SI_EQ_1, NOTIFIER);
     $width(negedge CDN &&& D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$CDN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(posedge CP &&& CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwh$CP$CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(negedge CP &&& CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$CP$CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_SDF03D1 (Q, QN, CP, D, SDN, SE, SI);
input  CP ;
input  D ;
input  SDN ;
input  SE ;
input  SI ;
output Q ;
output QN ;
reg NOTIFIER ;
reg ReSeT;

`ifdef  RSTn_lib
	 initial begin
		ReSeT = 0 ;
		#3 ReSeT = 1 ;
		#111 ReSeT = 0 ;
	end
  `else initial  ReSeT = 0;
`endif

   udp_mux2 (I0_D, D, SI, SE);
   not (I0_SET, SDN);
   udp_dff (N_S_XM29_G, I0_D, CP, ReSeT/*1'B0*/, I0_SET, NOTIFIER);
   not (N_NET0130_XM26_D, N_S_XM29_G);
   buf (Q, N_S_XM29_G);
   not (QN, N_S_XM29_G);
   and (SDN_EQ_1_AN_SE_EQ_1, SDN, SE);
   not (I9_out, D);
   not (I10_out, SE);
   not (I12_out, SI);
   and (D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, I9_out, I10_out, I12_out);
   not (I14_out, SE);
   and (SDN_EQ_1_AN_SE_EQ_0, SDN, I14_out);
   not (I16_out, D);
   not (I18_out, SE);
   not (I20_out, SI);
   and (D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, I16_out, SDN, I18_out, I20_out);

   specify
     // delay parameters
     specparam
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tpllh$CP$QN = 1.0,
       tplhl$CP$QN = 1.0,
       tphlh$SDN$Q = 1.0,
       tphhl$SDN$QN = 1.0,
       tminpwh$CP$D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwl$CP$D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwl$SDN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tsetup_negedge$D$CP$SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       thold_negedge$D$CP$SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       tsetup_negedge$SE$CP$SDN_EQ_1 = 1.0,
       thold_negedge$SE$CP$SDN_EQ_1 = 1.0,
       tsetup_negedge$SI$CP$SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       thold_negedge$SI$CP$SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       tsetup_posedge$D$CP$SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       thold_posedge$D$CP$SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       tsetup_posedge$SE$CP$SDN_EQ_1 = 1.0,
       thold_posedge$SE$CP$SDN_EQ_1 = 1.0,
       tsetup_posedge$SI$CP$SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       thold_posedge$SI$CP$SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       trec$SDN$CP$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       trem$SDN$CP$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0;

     // path delays
     (posedge CP *> (QN -: SE?SI:D)) = (tpllh$CP$QN, tplhl$CP$QN);
     (posedge CP *> (Q +: SE?SI:D)) = (tpllh$CP$Q, tplhl$CP$Q);
     (negedge SDN *> (QN -: 1'b1)) = (0, tphhl$SDN$QN);
     (negedge SDN *> (Q +: 1'b1)) = (tphlh$SDN$Q, 0);
     $setuphold(posedge CP &&& SDN_EQ_1_AN_SE_EQ_0 == 1'b1, negedge D, tsetup_negedge$D$CP$SDN_EQ_1_AN_SE_EQ_0, thold_negedge$D$CP$SDN_EQ_1_AN_SE_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& SDN == 1'b1, negedge SE, tsetup_negedge$SE$CP$SDN_EQ_1, thold_negedge$SE$CP$SDN_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& SDN_EQ_1_AN_SE_EQ_1 == 1'b1, negedge SI, tsetup_negedge$SI$CP$SDN_EQ_1_AN_SE_EQ_1, thold_negedge$SI$CP$SDN_EQ_1_AN_SE_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& SDN_EQ_1_AN_SE_EQ_0 == 1'b1, posedge D, tsetup_posedge$D$CP$SDN_EQ_1_AN_SE_EQ_0, thold_posedge$D$CP$SDN_EQ_1_AN_SE_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& SDN == 1'b1, posedge SE, tsetup_posedge$SE$CP$SDN_EQ_1, thold_posedge$SE$CP$SDN_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& SDN_EQ_1_AN_SE_EQ_1 == 1'b1, posedge SI, tsetup_posedge$SI$CP$SDN_EQ_1_AN_SE_EQ_1, thold_posedge$SI$CP$SDN_EQ_1_AN_SE_EQ_1, NOTIFIER);
     $recrem(posedge SDN, posedge CP &&& D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, trec$SDN$CP$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, trem$SDN$CP$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, NOTIFIER);
     $width(posedge CP &&& D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwh$CP$D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(negedge CP &&& D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$CP$D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(negedge SDN &&& D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$SDN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_SDF03D2 (Q, QN, CP, D, SDN, SE, SI);
input  CP ;
input  D ;
input  SDN ;
input  SE ;
input  SI ;
output Q ;
output QN ;
reg NOTIFIER ;

   udp_mux2 (I0_D, D, SI, SE);
   not (I0_SET, SDN);
   udp_dff (N_S_XM29_G, I0_D, CP, 1'B0, I0_SET, NOTIFIER);
   not (N_NET0130_XM26_D, N_S_XM29_G);
   buf (Q, N_S_XM29_G);
   not (QN, N_S_XM29_G);
   and (SDN_EQ_1_AN_SE_EQ_1, SDN, SE);
   not (I9_out, D);
   not (I10_out, SE);
   not (I12_out, SI);
   and (D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, I9_out, I10_out, I12_out);
   not (I14_out, SE);
   and (SDN_EQ_1_AN_SE_EQ_0, SDN, I14_out);
   not (I16_out, D);
   not (I18_out, SE);
   not (I20_out, SI);
   and (D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, I16_out, SDN, I18_out, I20_out);

   specify
     // delay parameters
     specparam
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tpllh$CP$QN = 1.0,
       tplhl$CP$QN = 1.0,
       tphlh$SDN$Q = 1.0,
       tphhl$SDN$QN = 1.0,
       tminpwh$CP$D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwl$CP$D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwl$SDN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tsetup_negedge$D$CP$SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       thold_negedge$D$CP$SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       tsetup_negedge$SE$CP$SDN_EQ_1 = 1.0,
       thold_negedge$SE$CP$SDN_EQ_1 = 1.0,
       tsetup_negedge$SI$CP$SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       thold_negedge$SI$CP$SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       tsetup_posedge$D$CP$SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       thold_posedge$D$CP$SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       tsetup_posedge$SE$CP$SDN_EQ_1 = 1.0,
       thold_posedge$SE$CP$SDN_EQ_1 = 1.0,
       tsetup_posedge$SI$CP$SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       thold_posedge$SI$CP$SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       trec$SDN$CP$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       trem$SDN$CP$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0;

     // path delays
     (posedge CP *> (QN -: SE?SI:D)) = (tpllh$CP$QN, tplhl$CP$QN);
     (posedge CP *> (Q +: SE?SI:D)) = (tpllh$CP$Q, tplhl$CP$Q);
     (negedge SDN *> (QN -: 1'b1)) = (0, tphhl$SDN$QN);
     (negedge SDN *> (Q +: 1'b1)) = (tphlh$SDN$Q, 0);
     $setuphold(posedge CP &&& SDN_EQ_1_AN_SE_EQ_0 == 1'b1, negedge D, tsetup_negedge$D$CP$SDN_EQ_1_AN_SE_EQ_0, thold_negedge$D$CP$SDN_EQ_1_AN_SE_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& SDN == 1'b1, negedge SE, tsetup_negedge$SE$CP$SDN_EQ_1, thold_negedge$SE$CP$SDN_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& SDN_EQ_1_AN_SE_EQ_1 == 1'b1, negedge SI, tsetup_negedge$SI$CP$SDN_EQ_1_AN_SE_EQ_1, thold_negedge$SI$CP$SDN_EQ_1_AN_SE_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& SDN_EQ_1_AN_SE_EQ_0 == 1'b1, posedge D, tsetup_posedge$D$CP$SDN_EQ_1_AN_SE_EQ_0, thold_posedge$D$CP$SDN_EQ_1_AN_SE_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& SDN == 1'b1, posedge SE, tsetup_posedge$SE$CP$SDN_EQ_1, thold_posedge$SE$CP$SDN_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& SDN_EQ_1_AN_SE_EQ_1 == 1'b1, posedge SI, tsetup_posedge$SI$CP$SDN_EQ_1_AN_SE_EQ_1, thold_posedge$SI$CP$SDN_EQ_1_AN_SE_EQ_1, NOTIFIER);
     $recrem(posedge SDN, posedge CP &&& D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, trec$SDN$CP$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, trem$SDN$CP$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, NOTIFIER);
     $width(posedge CP &&& D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwh$CP$D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(negedge CP &&& D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$CP$D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(negedge SDN &&& D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$SDN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_SDF03D4 (Q, QN, CP, D, SDN, SE, SI);
input  CP ;
input  D ;
input  SDN ;
input  SE ;
input  SI ;
output Q ;
output QN ;
reg NOTIFIER ;

   udp_mux2 (I0_D, D, SI, SE);
   not (I0_SET, SDN);
   udp_dff (N_S_XM29_G, I0_D, CP, 1'B0, I0_SET, NOTIFIER);
   not (N_NET0130_XM26_D, N_S_XM29_G);
   buf (Q, N_S_XM29_G);
   not (QN, N_S_XM29_G);
   and (SDN_EQ_1_AN_SE_EQ_1, SDN, SE);
   not (I9_out, D);
   not (I10_out, SE);
   not (I12_out, SI);
   and (D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, I9_out, I10_out, I12_out);
   not (I14_out, SE);
   and (SDN_EQ_1_AN_SE_EQ_0, SDN, I14_out);
   not (I16_out, D);
   not (I18_out, SE);
   not (I20_out, SI);
   and (D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, I16_out, SDN, I18_out, I20_out);

   specify
     // delay parameters
     specparam
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tpllh$CP$QN = 1.0,
       tplhl$CP$QN = 1.0,
       tphlh$SDN$Q = 1.0,
       tphhl$SDN$QN = 1.0,
       tminpwh$CP$D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwl$CP$D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwl$SDN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tsetup_negedge$D$CP$SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       thold_negedge$D$CP$SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       tsetup_negedge$SE$CP$SDN_EQ_1 = 1.0,
       thold_negedge$SE$CP$SDN_EQ_1 = 1.0,
       tsetup_negedge$SI$CP$SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       thold_negedge$SI$CP$SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       tsetup_posedge$D$CP$SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       thold_posedge$D$CP$SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       tsetup_posedge$SE$CP$SDN_EQ_1 = 1.0,
       thold_posedge$SE$CP$SDN_EQ_1 = 1.0,
       tsetup_posedge$SI$CP$SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       thold_posedge$SI$CP$SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       trec$SDN$CP$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       trem$SDN$CP$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0;

     // path delays
     (posedge CP *> (QN -: SE?SI:D)) = (tpllh$CP$QN, tplhl$CP$QN);
     (posedge CP *> (Q +: SE?SI:D)) = (tpllh$CP$Q, tplhl$CP$Q);
     (negedge SDN *> (QN -: 1'b1)) = (0, tphhl$SDN$QN);
     (negedge SDN *> (Q +: 1'b1)) = (tphlh$SDN$Q, 0);
     $setuphold(posedge CP &&& SDN_EQ_1_AN_SE_EQ_0 == 1'b1, negedge D, tsetup_negedge$D$CP$SDN_EQ_1_AN_SE_EQ_0, thold_negedge$D$CP$SDN_EQ_1_AN_SE_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& SDN == 1'b1, negedge SE, tsetup_negedge$SE$CP$SDN_EQ_1, thold_negedge$SE$CP$SDN_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& SDN_EQ_1_AN_SE_EQ_1 == 1'b1, negedge SI, tsetup_negedge$SI$CP$SDN_EQ_1_AN_SE_EQ_1, thold_negedge$SI$CP$SDN_EQ_1_AN_SE_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& SDN_EQ_1_AN_SE_EQ_0 == 1'b1, posedge D, tsetup_posedge$D$CP$SDN_EQ_1_AN_SE_EQ_0, thold_posedge$D$CP$SDN_EQ_1_AN_SE_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& SDN == 1'b1, posedge SE, tsetup_posedge$SE$CP$SDN_EQ_1, thold_posedge$SE$CP$SDN_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& SDN_EQ_1_AN_SE_EQ_1 == 1'b1, posedge SI, tsetup_posedge$SI$CP$SDN_EQ_1_AN_SE_EQ_1, thold_posedge$SI$CP$SDN_EQ_1_AN_SE_EQ_1, NOTIFIER);
     $recrem(posedge SDN, posedge CP &&& D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, trec$SDN$CP$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, trem$SDN$CP$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, NOTIFIER);
     $width(posedge CP &&& D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwh$CP$D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(negedge CP &&& D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$CP$D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(negedge SDN &&& D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$SDN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_SDF04D1 (Q, QN, CDN, CP, D, SDN, SE, SI);
input  CDN ;
input  CP ;
input  D ;
input  SDN ;
input  SE ;
input  SI ;
output Q ;
output QN ;
reg NOTIFIER ;

   udp_mux2 (I0_D, D, SI, SE);
   not (I0_CLEAR, CDN);
   not (I0_SET, SDN);
   udp_dff (N_S_XM33_G, I0_D, CP, I0_CLEAR, I0_SET, NOTIFIER);
   not (N_NET0130_XM30_D, N_S_XM33_G);
   not (Q, N_NET0130_XM30_D);
   buf (QN, N_NET0130_XM30_D);
   and (CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1, CDN, SDN, SE);
   and (CDN_EQ_1_AN_SDN_EQ_1, CDN, SDN);
   not (I13_out, SE);
   and (CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0, CDN, SDN, I13_out);
   not (I15_out, D);
   not (I16_out, SE);
   not (I18_out, SI);
   and (D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, I15_out, I16_out, I18_out);
   not (I20_out, D);
   not (I22_out, SE);
   not (I24_out, SI);
   and (D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, I20_out, SDN, I22_out, I24_out);
   not (I26_out, D);
   not (I29_out, SE);
   not (I31_out, SI);
   and (CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, CDN, I26_out, SDN, I29_out, I31_out);
   not (I33_out, CDN);
   not (I34_out, D);
   not (I36_out, SE);
   not (I38_out, SI);
   and (CDN_EQ_0_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, I33_out, I34_out, I36_out, I38_out);

   specify
     // delay parameters
     specparam
       tphhl$CDN$Q = 1.0,
       tphlh$CDN$QN = 1.0,
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tpllh$CP$QN = 1.0,
       tplhl$CP$QN = 1.0,
       tplhl$SDN$Q = 1.0,
       tphlh$SDN$Q = 1.0,
       tpllh$SDN$QN = 1.0,
       tphhl$SDN$QN = 1.0,
       tminpwl$CDN$D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwh$CP$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwl$CP$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwl$SDN$CDN_EQ_0_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tsetup_negedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       thold_negedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       tsetup_negedge$SE$CP$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       thold_negedge$SE$CP$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       tsetup_negedge$SI$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       thold_negedge$SI$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       tsetup_posedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       thold_posedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       tsetup_posedge$SE$CP$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       thold_posedge$SE$CP$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       tsetup_posedge$SI$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       thold_posedge$SI$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       trec$CDN$CP$SDN_EQ_1 = 1.0,
       trem$CDN$CP$SDN_EQ_1 = 1.0,
       trec$CDN$SDN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       trec$SDN$CP$CDN_EQ_1 = 1.0,
       trem$SDN$CP$CDN_EQ_1 = 1.0;

     // path delays
     (posedge CP *> (QN -: SE?SI:D)) = (tpllh$CP$QN, tplhl$CP$QN);
     (posedge CP *> (Q +: SE?SI:D)) = (tpllh$CP$Q, tplhl$CP$Q);
     (negedge SDN *> (QN -: 1'b1)) = (tpllh$SDN$QN, tphhl$SDN$QN);
     (negedge SDN *> (Q +: 1'b1)) = (tphlh$SDN$Q, tplhl$SDN$Q);
     (negedge CDN *> (QN +: 1'b1)) = (tphlh$CDN$QN, 0);
     (negedge CDN *> (Q -: 1'b1)) = (0, tphhl$CDN$Q);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0 == 1'b1, negedge D, tsetup_negedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0, thold_negedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_SDN_EQ_1 == 1'b1, negedge SE, tsetup_negedge$SE$CP$CDN_EQ_1_AN_SDN_EQ_1, thold_negedge$SE$CP$CDN_EQ_1_AN_SDN_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1 == 1'b1, negedge SI, tsetup_negedge$SI$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1, thold_negedge$SI$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0 == 1'b1, posedge D, tsetup_posedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0, thold_posedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_SDN_EQ_1 == 1'b1, posedge SE, tsetup_posedge$SE$CP$CDN_EQ_1_AN_SDN_EQ_1, thold_posedge$SE$CP$CDN_EQ_1_AN_SDN_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1 == 1'b1, posedge SI, tsetup_posedge$SI$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1, thold_posedge$SI$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1, NOTIFIER);
     $recrem(posedge CDN, posedge CP &&& SDN == 1'b1, trec$CDN$CP$SDN_EQ_1, trem$CDN$CP$SDN_EQ_1, NOTIFIER);
     $recovery(posedge CDN, posedge SDN &&& D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, trec$CDN$SDN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, NOTIFIER);
     $recrem(posedge SDN, posedge CP &&& CDN == 1'b1, trec$SDN$CP$CDN_EQ_1, trem$SDN$CP$CDN_EQ_1, NOTIFIER);
     $width(negedge CDN &&& D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$CDN$D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(posedge CP &&& CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwh$CP$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(negedge CP &&& CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$CP$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(negedge SDN &&& CDN_EQ_0_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$SDN$CDN_EQ_0_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_SDF04D2 (Q, QN, CDN, CP, D, SDN, SE, SI);
input  CDN ;
input  CP ;
input  D ;
input  SDN ;
input  SE ;
input  SI ;
output Q ;
output QN ;
reg NOTIFIER ;

   udp_mux2 (I0_D, D, SI, SE);
   not (I0_CLEAR, CDN);
   not (I0_SET, SDN);
   udp_dff (N_S_XM33_G, I0_D, CP, I0_CLEAR, I0_SET, NOTIFIER);
   not (N_NET0130_XM30_D, N_S_XM33_G);
   not (Q, N_NET0130_XM30_D);
   buf (QN, N_NET0130_XM30_D);
   and (CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1, CDN, SDN, SE);
   and (CDN_EQ_1_AN_SDN_EQ_1, CDN, SDN);
   not (I13_out, SE);
   and (CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0, CDN, SDN, I13_out);
   not (I15_out, D);
   not (I16_out, SE);
   not (I18_out, SI);
   and (D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, I15_out, I16_out, I18_out);
   not (I20_out, D);
   not (I22_out, SE);
   not (I24_out, SI);
   and (D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, I20_out, SDN, I22_out, I24_out);
   not (I26_out, D);
   not (I29_out, SE);
   not (I31_out, SI);
   and (CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, CDN, I26_out, SDN, I29_out, I31_out);
   not (I33_out, CDN);
   not (I34_out, D);
   not (I36_out, SE);
   not (I38_out, SI);
   and (CDN_EQ_0_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, I33_out, I34_out, I36_out, I38_out);

   specify
     // delay parameters
     specparam
       tphhl$CDN$Q = 1.0,
       tphlh$CDN$QN = 1.0,
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tpllh$CP$QN = 1.0,
       tplhl$CP$QN = 1.0,
       tplhl$SDN$Q = 1.0,
       tphlh$SDN$Q = 1.0,
       tpllh$SDN$QN = 1.0,
       tphhl$SDN$QN = 1.0,
       tminpwl$CDN$D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwh$CP$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwl$CP$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwl$SDN$CDN_EQ_0_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tsetup_negedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       thold_negedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       tsetup_negedge$SE$CP$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       thold_negedge$SE$CP$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       tsetup_negedge$SI$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       thold_negedge$SI$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       tsetup_posedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       thold_posedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       tsetup_posedge$SE$CP$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       thold_posedge$SE$CP$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       tsetup_posedge$SI$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       thold_posedge$SI$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       trec$CDN$CP$SDN_EQ_1 = 1.0,
       trem$CDN$CP$SDN_EQ_1 = 1.0,
       trec$CDN$SDN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       trec$SDN$CP$CDN_EQ_1 = 1.0,
       trem$SDN$CP$CDN_EQ_1 = 1.0;

     // path delays
     (posedge CP *> (QN -: SE?SI:D)) = (tpllh$CP$QN, tplhl$CP$QN);
     (posedge CP *> (Q +: SE?SI:D)) = (tpllh$CP$Q, tplhl$CP$Q);
     (negedge SDN *> (QN -: 1'b1)) = (tpllh$SDN$QN, tphhl$SDN$QN);
     (negedge SDN *> (Q +: 1'b1)) = (tphlh$SDN$Q, tplhl$SDN$Q);
     (negedge CDN *> (QN +: 1'b1)) = (tphlh$CDN$QN, 0);
     (negedge CDN *> (Q -: 1'b1)) = (0, tphhl$CDN$Q);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0 == 1'b1, negedge D, tsetup_negedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0, thold_negedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_SDN_EQ_1 == 1'b1, negedge SE, tsetup_negedge$SE$CP$CDN_EQ_1_AN_SDN_EQ_1, thold_negedge$SE$CP$CDN_EQ_1_AN_SDN_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1 == 1'b1, negedge SI, tsetup_negedge$SI$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1, thold_negedge$SI$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0 == 1'b1, posedge D, tsetup_posedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0, thold_posedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_SDN_EQ_1 == 1'b1, posedge SE, tsetup_posedge$SE$CP$CDN_EQ_1_AN_SDN_EQ_1, thold_posedge$SE$CP$CDN_EQ_1_AN_SDN_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1 == 1'b1, posedge SI, tsetup_posedge$SI$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1, thold_posedge$SI$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1, NOTIFIER);
     $recrem(posedge CDN, posedge CP &&& SDN == 1'b1, trec$CDN$CP$SDN_EQ_1, trem$CDN$CP$SDN_EQ_1, NOTIFIER);
     $recovery(posedge CDN, posedge SDN &&& D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, trec$CDN$SDN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, NOTIFIER);
     $recrem(posedge SDN, posedge CP &&& CDN == 1'b1, trec$SDN$CP$CDN_EQ_1, trem$SDN$CP$CDN_EQ_1, NOTIFIER);
     $width(negedge CDN &&& D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$CDN$D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(posedge CP &&& CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwh$CP$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(negedge CP &&& CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$CP$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(negedge SDN &&& CDN_EQ_0_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$SDN$CDN_EQ_0_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_SDF04D4 (Q, QN, CDN, CP, D, SDN, SE, SI);
input  CDN ;
input  CP ;
input  D ;
input  SDN ;
input  SE ;
input  SI ;
output Q ;
output QN ;
reg NOTIFIER ;

   udp_mux2 (I0_D, D, SI, SE);
   not (I0_CLEAR, CDN);
   not (I0_SET, SDN);
   udp_dff (N_S_XM33_G, I0_D, CP, I0_CLEAR, I0_SET, NOTIFIER);
   not (N_NET0130_XM30_D, N_S_XM33_G);
   not (Q, N_NET0130_XM30_D);
   buf (QN, N_NET0130_XM30_D);
   and (CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1, CDN, SDN, SE);
   and (CDN_EQ_1_AN_SDN_EQ_1, CDN, SDN);
   not (I13_out, SE);
   and (CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0, CDN, SDN, I13_out);
   not (I15_out, D);
   not (I16_out, SE);
   not (I18_out, SI);
   and (D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, I15_out, I16_out, I18_out);
   not (I20_out, D);
   not (I22_out, SE);
   not (I24_out, SI);
   and (D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, I20_out, SDN, I22_out, I24_out);
   not (I26_out, D);
   not (I29_out, SE);
   not (I31_out, SI);
   and (CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, CDN, I26_out, SDN, I29_out, I31_out);
   not (I33_out, CDN);
   not (I34_out, D);
   not (I36_out, SE);
   not (I38_out, SI);
   and (CDN_EQ_0_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, I33_out, I34_out, I36_out, I38_out);

   specify
     // delay parameters
     specparam
       tphhl$CDN$Q = 1.0,
       tphlh$CDN$QN = 1.0,
       tpllh$CP$Q = 1.0,
       tplhl$CP$Q = 1.0,
       tpllh$CP$QN = 1.0,
       tplhl$CP$QN = 1.0,
       tplhl$SDN$Q = 1.0,
       tphlh$SDN$Q = 1.0,
       tpllh$SDN$QN = 1.0,
       tphhl$SDN$QN = 1.0,
       tminpwl$CDN$D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwh$CP$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwl$CP$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwl$SDN$CDN_EQ_0_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tsetup_negedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       thold_negedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       tsetup_negedge$SE$CP$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       thold_negedge$SE$CP$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       tsetup_negedge$SI$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       thold_negedge$SI$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       tsetup_posedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       thold_posedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       tsetup_posedge$SE$CP$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       thold_posedge$SE$CP$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       tsetup_posedge$SI$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       thold_posedge$SI$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       trec$CDN$CP$SDN_EQ_1 = 1.0,
       trem$CDN$CP$SDN_EQ_1 = 1.0,
       trec$CDN$SDN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       trec$SDN$CP$CDN_EQ_1 = 1.0,
       trem$SDN$CP$CDN_EQ_1 = 1.0;

     // path delays
     (posedge CP *> (QN -: SE?SI:D)) = (tpllh$CP$QN, tplhl$CP$QN);
     (posedge CP *> (Q +: SE?SI:D)) = (tpllh$CP$Q, tplhl$CP$Q);
     (negedge SDN *> (QN -: 1'b1)) = (tpllh$SDN$QN, tphhl$SDN$QN);
     (negedge SDN *> (Q +: 1'b1)) = (tphlh$SDN$Q, tplhl$SDN$Q);
     (negedge CDN *> (QN +: 1'b1)) = (tphlh$CDN$QN, 0);
     (negedge CDN *> (Q -: 1'b1)) = (0, tphhl$CDN$Q);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0 == 1'b1, negedge D, tsetup_negedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0, thold_negedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_SDN_EQ_1 == 1'b1, negedge SE, tsetup_negedge$SE$CP$CDN_EQ_1_AN_SDN_EQ_1, thold_negedge$SE$CP$CDN_EQ_1_AN_SDN_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1 == 1'b1, negedge SI, tsetup_negedge$SI$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1, thold_negedge$SI$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0 == 1'b1, posedge D, tsetup_posedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0, thold_posedge$D$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0, NOTIFIER);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_SDN_EQ_1 == 1'b1, posedge SE, tsetup_posedge$SE$CP$CDN_EQ_1_AN_SDN_EQ_1, thold_posedge$SE$CP$CDN_EQ_1_AN_SDN_EQ_1, NOTIFIER);
     $setuphold(posedge CP &&& CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1 == 1'b1, posedge SI, tsetup_posedge$SI$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1, thold_posedge$SI$CP$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1, NOTIFIER);
     $recrem(posedge CDN, posedge CP &&& SDN == 1'b1, trec$CDN$CP$SDN_EQ_1, trem$CDN$CP$SDN_EQ_1, NOTIFIER);
     $recovery(posedge CDN, posedge SDN &&& D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, trec$CDN$SDN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, NOTIFIER);
     $recrem(posedge SDN, posedge CP &&& CDN == 1'b1, trec$SDN$CP$CDN_EQ_1, trem$SDN$CP$CDN_EQ_1, NOTIFIER);
     $width(negedge CDN &&& D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$CDN$D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(posedge CP &&& CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwh$CP$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(negedge CP &&& CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$CP$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(negedge SDN &&& CDN_EQ_0_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$SDN$CDN_EQ_0_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_SDF05D1 (Q, QN, CPN, D, SE, SI);
input  CPN ;
input  D ;
input  SE ;
input  SI ;
output Q ;
output QN ;
reg NOTIFIER ;

   udp_mux2 (I0_D, D, SI, SE);
   not (I0_CLOCK, CPN);
   udp_dff (N_S_XM27_G, I0_D, I0_CLOCK, 1'B0, 1'B0, NOTIFIER);
   not (N_NET0130_XM24_D, N_S_XM27_G);
   buf (Q, N_S_XM27_G);
   not (QN, N_S_XM27_G);
   not (I8_out, D);
   and (D_EQ_0_AN_SI_EQ_1, I8_out, SI);
   not (I10_out, SI);
   and (D_EQ_1_AN_SI_EQ_0, D, I10_out);
   not (I12_out, D);
   not (I13_out, SE);
   not (I15_out, SI);
   and (D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, I12_out, I13_out, I15_out);

   specify
     // delay parameters
     specparam
       tphlh$CPN$Q = 1.0,
       tphhl$CPN$Q = 1.0,
       tphlh$CPN$QN = 1.0,
       tphhl$CPN$QN = 1.0,
       tminpwh$CPN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwl$CPN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tsetup_negedge$D$CPN$SE_EQ_0 = 1.0,
       thold_negedge$D$CPN$SE_EQ_0 = 1.0,
       tsetup_negedge$SE$CPN$D_EQ_0_AN_SI_EQ_1 = 1.0,
       thold_negedge$SE$CPN$D_EQ_0_AN_SI_EQ_1 = 1.0,
       tsetup_negedge$SE$CPN$D_EQ_1_AN_SI_EQ_0 = 1.0,
       thold_negedge$SE$CPN$D_EQ_1_AN_SI_EQ_0 = 1.0,
       tsetup_negedge$SI$CPN$SE_EQ_1 = 1.0,
       thold_negedge$SI$CPN$SE_EQ_1 = 1.0,
       tsetup_posedge$D$CPN$SE_EQ_0 = 1.0,
       thold_posedge$D$CPN$SE_EQ_0 = 1.0,
       tsetup_posedge$SE$CPN$D_EQ_0_AN_SI_EQ_1 = 1.0,
       thold_posedge$SE$CPN$D_EQ_0_AN_SI_EQ_1 = 1.0,
       tsetup_posedge$SE$CPN$D_EQ_1_AN_SI_EQ_0 = 1.0,
       thold_posedge$SE$CPN$D_EQ_1_AN_SI_EQ_0 = 1.0,
       tsetup_posedge$SI$CPN$SE_EQ_1 = 1.0,
       thold_posedge$SI$CPN$SE_EQ_1 = 1.0;

     // path delays
     (negedge CPN *> (QN -: SE?SI:D)) = (tphlh$CPN$QN, tphhl$CPN$QN);
     (negedge CPN *> (Q +: SE?SI:D)) = (tphlh$CPN$Q, tphhl$CPN$Q);
     $setuphold(negedge CPN &&& SE == 1'b0, negedge D, tsetup_negedge$D$CPN$SE_EQ_0, thold_negedge$D$CPN$SE_EQ_0, NOTIFIER);
     $setuphold(negedge CPN &&& D_EQ_0_AN_SI_EQ_1 == 1'b1, negedge SE, tsetup_negedge$SE$CPN$D_EQ_0_AN_SI_EQ_1, thold_negedge$SE$CPN$D_EQ_0_AN_SI_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& D_EQ_1_AN_SI_EQ_0 == 1'b1, negedge SE, tsetup_negedge$SE$CPN$D_EQ_1_AN_SI_EQ_0, thold_negedge$SE$CPN$D_EQ_1_AN_SI_EQ_0, NOTIFIER);
     $setuphold(negedge CPN &&& SE == 1'b1, negedge SI, tsetup_negedge$SI$CPN$SE_EQ_1, thold_negedge$SI$CPN$SE_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& SE == 1'b0, posedge D, tsetup_posedge$D$CPN$SE_EQ_0, thold_posedge$D$CPN$SE_EQ_0, NOTIFIER);
     $setuphold(negedge CPN &&& D_EQ_0_AN_SI_EQ_1 == 1'b1, posedge SE, tsetup_posedge$SE$CPN$D_EQ_0_AN_SI_EQ_1, thold_posedge$SE$CPN$D_EQ_0_AN_SI_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& D_EQ_1_AN_SI_EQ_0 == 1'b1, posedge SE, tsetup_posedge$SE$CPN$D_EQ_1_AN_SI_EQ_0, thold_posedge$SE$CPN$D_EQ_1_AN_SI_EQ_0, NOTIFIER);
     $setuphold(negedge CPN &&& SE == 1'b1, posedge SI, tsetup_posedge$SI$CPN$SE_EQ_1, thold_posedge$SI$CPN$SE_EQ_1, NOTIFIER);
     $width(posedge CPN &&& D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwh$CPN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(negedge CPN &&& D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$CPN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_SDF05D2 (Q, QN, CPN, D, SE, SI);
input  CPN ;
input  D ;
input  SE ;
input  SI ;
output Q ;
output QN ;
reg NOTIFIER ;

   udp_mux2 (I0_D, D, SI, SE);
   not (I0_CLOCK, CPN);
   udp_dff (N_S_XM27_G, I0_D, I0_CLOCK, 1'B0, 1'B0, NOTIFIER);
   not (N_NET0130_XM24_D, N_S_XM27_G);
   buf (Q, N_S_XM27_G);
   not (QN, N_S_XM27_G);
   not (I8_out, D);
   and (D_EQ_0_AN_SI_EQ_1, I8_out, SI);
   not (I10_out, SI);
   and (D_EQ_1_AN_SI_EQ_0, D, I10_out);
   not (I12_out, D);
   not (I13_out, SE);
   not (I15_out, SI);
   and (D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, I12_out, I13_out, I15_out);

   specify
     // delay parameters
     specparam
       tphlh$CPN$Q = 1.0,
       tphhl$CPN$Q = 1.0,
       tphlh$CPN$QN = 1.0,
       tphhl$CPN$QN = 1.0,
       tminpwh$CPN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwl$CPN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tsetup_negedge$D$CPN$SE_EQ_0 = 1.0,
       thold_negedge$D$CPN$SE_EQ_0 = 1.0,
       tsetup_negedge$SE$CPN$D_EQ_0_AN_SI_EQ_1 = 1.0,
       thold_negedge$SE$CPN$D_EQ_0_AN_SI_EQ_1 = 1.0,
       tsetup_negedge$SE$CPN$D_EQ_1_AN_SI_EQ_0 = 1.0,
       thold_negedge$SE$CPN$D_EQ_1_AN_SI_EQ_0 = 1.0,
       tsetup_negedge$SI$CPN$SE_EQ_1 = 1.0,
       thold_negedge$SI$CPN$SE_EQ_1 = 1.0,
       tsetup_posedge$D$CPN$SE_EQ_0 = 1.0,
       thold_posedge$D$CPN$SE_EQ_0 = 1.0,
       tsetup_posedge$SE$CPN$D_EQ_0_AN_SI_EQ_1 = 1.0,
       thold_posedge$SE$CPN$D_EQ_0_AN_SI_EQ_1 = 1.0,
       tsetup_posedge$SE$CPN$D_EQ_1_AN_SI_EQ_0 = 1.0,
       thold_posedge$SE$CPN$D_EQ_1_AN_SI_EQ_0 = 1.0,
       tsetup_posedge$SI$CPN$SE_EQ_1 = 1.0,
       thold_posedge$SI$CPN$SE_EQ_1 = 1.0;

     // path delays
     (negedge CPN *> (QN -: SE?SI:D)) = (tphlh$CPN$QN, tphhl$CPN$QN);
     (negedge CPN *> (Q +: SE?SI:D)) = (tphlh$CPN$Q, tphhl$CPN$Q);
     $setuphold(negedge CPN &&& SE == 1'b0, negedge D, tsetup_negedge$D$CPN$SE_EQ_0, thold_negedge$D$CPN$SE_EQ_0, NOTIFIER);
     $setuphold(negedge CPN &&& D_EQ_0_AN_SI_EQ_1 == 1'b1, negedge SE, tsetup_negedge$SE$CPN$D_EQ_0_AN_SI_EQ_1, thold_negedge$SE$CPN$D_EQ_0_AN_SI_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& D_EQ_1_AN_SI_EQ_0 == 1'b1, negedge SE, tsetup_negedge$SE$CPN$D_EQ_1_AN_SI_EQ_0, thold_negedge$SE$CPN$D_EQ_1_AN_SI_EQ_0, NOTIFIER);
     $setuphold(negedge CPN &&& SE == 1'b1, negedge SI, tsetup_negedge$SI$CPN$SE_EQ_1, thold_negedge$SI$CPN$SE_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& SE == 1'b0, posedge D, tsetup_posedge$D$CPN$SE_EQ_0, thold_posedge$D$CPN$SE_EQ_0, NOTIFIER);
     $setuphold(negedge CPN &&& D_EQ_0_AN_SI_EQ_1 == 1'b1, posedge SE, tsetup_posedge$SE$CPN$D_EQ_0_AN_SI_EQ_1, thold_posedge$SE$CPN$D_EQ_0_AN_SI_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& D_EQ_1_AN_SI_EQ_0 == 1'b1, posedge SE, tsetup_posedge$SE$CPN$D_EQ_1_AN_SI_EQ_0, thold_posedge$SE$CPN$D_EQ_1_AN_SI_EQ_0, NOTIFIER);
     $setuphold(negedge CPN &&& SE == 1'b1, posedge SI, tsetup_posedge$SI$CPN$SE_EQ_1, thold_posedge$SI$CPN$SE_EQ_1, NOTIFIER);
     $width(posedge CPN &&& D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwh$CPN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(negedge CPN &&& D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$CPN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_SDF05D4 (Q, QN, CPN, D, SE, SI);
input  CPN ;
input  D ;
input  SE ;
input  SI ;
output Q ;
output QN ;
reg NOTIFIER ;

   udp_mux2 (I0_D, D, SI, SE);
   not (I0_CLOCK, CPN);
   udp_dff (N_S_XM27_G, I0_D, I0_CLOCK, 1'B0, 1'B0, NOTIFIER);
   not (N_NET0130_XM24_D, N_S_XM27_G);
   buf (Q, N_S_XM27_G);
   not (QN, N_S_XM27_G);
   not (I8_out, D);
   and (D_EQ_0_AN_SI_EQ_1, I8_out, SI);
   not (I10_out, SI);
   and (D_EQ_1_AN_SI_EQ_0, D, I10_out);
   not (I12_out, D);
   not (I13_out, SE);
   not (I15_out, SI);
   and (D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, I12_out, I13_out, I15_out);

   specify
     // delay parameters
     specparam
       tphlh$CPN$Q = 1.0,
       tphhl$CPN$Q = 1.0,
       tphlh$CPN$QN = 1.0,
       tphhl$CPN$QN = 1.0,
       tminpwh$CPN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwl$CPN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tsetup_negedge$D$CPN$SE_EQ_0 = 1.0,
       thold_negedge$D$CPN$SE_EQ_0 = 1.0,
       tsetup_negedge$SE$CPN$D_EQ_0_AN_SI_EQ_1 = 1.0,
       thold_negedge$SE$CPN$D_EQ_0_AN_SI_EQ_1 = 1.0,
       tsetup_negedge$SE$CPN$D_EQ_1_AN_SI_EQ_0 = 1.0,
       thold_negedge$SE$CPN$D_EQ_1_AN_SI_EQ_0 = 1.0,
       tsetup_negedge$SI$CPN$SE_EQ_1 = 1.0,
       thold_negedge$SI$CPN$SE_EQ_1 = 1.0,
       tsetup_posedge$D$CPN$SE_EQ_0 = 1.0,
       thold_posedge$D$CPN$SE_EQ_0 = 1.0,
       tsetup_posedge$SE$CPN$D_EQ_0_AN_SI_EQ_1 = 1.0,
       thold_posedge$SE$CPN$D_EQ_0_AN_SI_EQ_1 = 1.0,
       tsetup_posedge$SE$CPN$D_EQ_1_AN_SI_EQ_0 = 1.0,
       thold_posedge$SE$CPN$D_EQ_1_AN_SI_EQ_0 = 1.0,
       tsetup_posedge$SI$CPN$SE_EQ_1 = 1.0,
       thold_posedge$SI$CPN$SE_EQ_1 = 1.0;

     // path delays
     (negedge CPN *> (QN -: SE?SI:D)) = (tphlh$CPN$QN, tphhl$CPN$QN);
     (negedge CPN *> (Q +: SE?SI:D)) = (tphlh$CPN$Q, tphhl$CPN$Q);
     $setuphold(negedge CPN &&& SE == 1'b0, negedge D, tsetup_negedge$D$CPN$SE_EQ_0, thold_negedge$D$CPN$SE_EQ_0, NOTIFIER);
     $setuphold(negedge CPN &&& D_EQ_0_AN_SI_EQ_1 == 1'b1, negedge SE, tsetup_negedge$SE$CPN$D_EQ_0_AN_SI_EQ_1, thold_negedge$SE$CPN$D_EQ_0_AN_SI_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& D_EQ_1_AN_SI_EQ_0 == 1'b1, negedge SE, tsetup_negedge$SE$CPN$D_EQ_1_AN_SI_EQ_0, thold_negedge$SE$CPN$D_EQ_1_AN_SI_EQ_0, NOTIFIER);
     $setuphold(negedge CPN &&& SE == 1'b1, negedge SI, tsetup_negedge$SI$CPN$SE_EQ_1, thold_negedge$SI$CPN$SE_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& SE == 1'b0, posedge D, tsetup_posedge$D$CPN$SE_EQ_0, thold_posedge$D$CPN$SE_EQ_0, NOTIFIER);
     $setuphold(negedge CPN &&& D_EQ_0_AN_SI_EQ_1 == 1'b1, posedge SE, tsetup_posedge$SE$CPN$D_EQ_0_AN_SI_EQ_1, thold_posedge$SE$CPN$D_EQ_0_AN_SI_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& D_EQ_1_AN_SI_EQ_0 == 1'b1, posedge SE, tsetup_posedge$SE$CPN$D_EQ_1_AN_SI_EQ_0, thold_posedge$SE$CPN$D_EQ_1_AN_SI_EQ_0, NOTIFIER);
     $setuphold(negedge CPN &&& SE == 1'b1, posedge SI, tsetup_posedge$SI$CPN$SE_EQ_1, thold_posedge$SI$CPN$SE_EQ_1, NOTIFIER);
     $width(posedge CPN &&& D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwh$CPN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(negedge CPN &&& D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$CPN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_SDF06D1 (Q, QN, CDN, CPN, D, SE, SI);
input  CDN ;
input  CPN ;
input  D ;
input  SE ;
input  SI ;
output Q ;
output QN ;
reg NOTIFIER ;

   udp_mux2 (I0_D, D, SI, SE);
   not (I0_CLOCK, CPN);
   not (I0_CLEAR, CDN);
   udp_dff (N_S_XM31_G, I0_D, I0_CLOCK, I0_CLEAR, 1'B0, NOTIFIER);
   not (N_NET0130_XM28_D, N_S_XM31_G);
   buf (Q, N_S_XM31_G);
   not (QN, N_S_XM31_G);
   and (CDN_EQ_1_AN_SE_EQ_1, CDN, SE);
   not (I10_out, SE);
   and (CDN_EQ_1_AN_SE_EQ_0, CDN, I10_out);
   not (I12_out, D);
   and (D_EQ_0_AN_SE_EQ_1_AN_SI_EQ_1, I12_out, SE, SI);
   not (I15_out, D);
   not (I16_out, SE);
   not (I18_out, SI);
   and (D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, I15_out, I16_out, I18_out);
   not (I20_out, D);
   not (I22_out, SE);
   not (I24_out, SI);
   and (CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, CDN, I20_out, I22_out, I24_out);

   specify
     // delay parameters
     specparam
       tphhl$CDN$Q = 1.0,
       tphlh$CDN$QN = 1.0,
       tphlh$CPN$Q = 1.0,
       tphhl$CPN$Q = 1.0,
       tphlh$CPN$QN = 1.0,
       tphhl$CPN$QN = 1.0,
       tminpwl$CDN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwh$CPN$CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwl$CPN$CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tsetup_negedge$D$CPN$CDN_EQ_1_AN_SE_EQ_0 = 1.0,
       thold_negedge$D$CPN$CDN_EQ_1_AN_SE_EQ_0 = 1.0,
       tsetup_negedge$SE$CPN$CDN_EQ_1 = 1.0,
       thold_negedge$SE$CPN$CDN_EQ_1 = 1.0,
       tsetup_negedge$SI$CPN$CDN_EQ_1_AN_SE_EQ_1 = 1.0,
       thold_negedge$SI$CPN$CDN_EQ_1_AN_SE_EQ_1 = 1.0,
       tsetup_posedge$D$CPN$CDN_EQ_1_AN_SE_EQ_0 = 1.0,
       thold_posedge$D$CPN$CDN_EQ_1_AN_SE_EQ_0 = 1.0,
       tsetup_posedge$SE$CPN$CDN_EQ_1 = 1.0,
       thold_posedge$SE$CPN$CDN_EQ_1 = 1.0,
       tsetup_posedge$SI$CPN$CDN_EQ_1_AN_SE_EQ_1 = 1.0,
       thold_posedge$SI$CPN$CDN_EQ_1_AN_SE_EQ_1 = 1.0,
       trec$CDN$CPN$D_EQ_0_AN_SE_EQ_1_AN_SI_EQ_1 = 1.0,
       trem$CDN$CPN$D_EQ_0_AN_SE_EQ_1_AN_SI_EQ_1 = 1.0;

     // path delays
     (negedge CPN *> (QN -: SE?SI:D)) = (tphlh$CPN$QN, tphhl$CPN$QN);
     (negedge CPN *> (Q +: SE?SI:D)) = (tphlh$CPN$Q, tphhl$CPN$Q);
     (negedge CDN *> (QN +: 1'b1)) = (tphlh$CDN$QN, 0);
     (negedge CDN *> (Q -: 1'b1)) = (0, tphhl$CDN$Q);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_SE_EQ_0 == 1'b1, negedge D, tsetup_negedge$D$CPN$CDN_EQ_1_AN_SE_EQ_0, thold_negedge$D$CPN$CDN_EQ_1_AN_SE_EQ_0, NOTIFIER);
     $setuphold(negedge CPN &&& CDN == 1'b1, negedge SE, tsetup_negedge$SE$CPN$CDN_EQ_1, thold_negedge$SE$CPN$CDN_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_SE_EQ_1 == 1'b1, negedge SI, tsetup_negedge$SI$CPN$CDN_EQ_1_AN_SE_EQ_1, thold_negedge$SI$CPN$CDN_EQ_1_AN_SE_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_SE_EQ_0 == 1'b1, posedge D, tsetup_posedge$D$CPN$CDN_EQ_1_AN_SE_EQ_0, thold_posedge$D$CPN$CDN_EQ_1_AN_SE_EQ_0, NOTIFIER);
     $setuphold(negedge CPN &&& CDN == 1'b1, posedge SE, tsetup_posedge$SE$CPN$CDN_EQ_1, thold_posedge$SE$CPN$CDN_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_SE_EQ_1 == 1'b1, posedge SI, tsetup_posedge$SI$CPN$CDN_EQ_1_AN_SE_EQ_1, thold_posedge$SI$CPN$CDN_EQ_1_AN_SE_EQ_1, NOTIFIER);
     $recrem(posedge CDN, negedge CPN &&& D_EQ_0_AN_SE_EQ_1_AN_SI_EQ_1 == 1'b1, trec$CDN$CPN$D_EQ_0_AN_SE_EQ_1_AN_SI_EQ_1, trem$CDN$CPN$D_EQ_0_AN_SE_EQ_1_AN_SI_EQ_1, NOTIFIER);
     $width(negedge CDN &&& D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$CDN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(posedge CPN &&& CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwh$CPN$CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(negedge CPN &&& CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$CPN$CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_SDF06D2 (Q, QN, CDN, CPN, D, SE, SI);
input  CDN ;
input  CPN ;
input  D ;
input  SE ;
input  SI ;
output Q ;
output QN ;
reg NOTIFIER ;

   udp_mux2 (I0_D, D, SI, SE);
   not (I0_CLOCK, CPN);
   not (I0_CLEAR, CDN);
   udp_dff (N_S_XM31_G, I0_D, I0_CLOCK, I0_CLEAR, 1'B0, NOTIFIER);
   not (N_NET0130_XM28_D, N_S_XM31_G);
   buf (Q, N_S_XM31_G);
   not (QN, N_S_XM31_G);
   and (CDN_EQ_1_AN_SE_EQ_1, CDN, SE);
   not (I10_out, SE);
   and (CDN_EQ_1_AN_SE_EQ_0, CDN, I10_out);
   not (I12_out, D);
   and (D_EQ_0_AN_SE_EQ_1_AN_SI_EQ_1, I12_out, SE, SI);
   not (I15_out, D);
   not (I16_out, SE);
   not (I18_out, SI);
   and (D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, I15_out, I16_out, I18_out);
   not (I20_out, D);
   not (I22_out, SE);
   not (I24_out, SI);
   and (CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, CDN, I20_out, I22_out, I24_out);

   specify
     // delay parameters
     specparam
       tphhl$CDN$Q = 1.0,
       tphlh$CDN$QN = 1.0,
       tphlh$CPN$Q = 1.0,
       tphhl$CPN$Q = 1.0,
       tphlh$CPN$QN = 1.0,
       tphhl$CPN$QN = 1.0,
       tminpwl$CDN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwh$CPN$CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwl$CPN$CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tsetup_negedge$D$CPN$CDN_EQ_1_AN_SE_EQ_0 = 1.0,
       thold_negedge$D$CPN$CDN_EQ_1_AN_SE_EQ_0 = 1.0,
       tsetup_negedge$SE$CPN$CDN_EQ_1 = 1.0,
       thold_negedge$SE$CPN$CDN_EQ_1 = 1.0,
       tsetup_negedge$SI$CPN$CDN_EQ_1_AN_SE_EQ_1 = 1.0,
       thold_negedge$SI$CPN$CDN_EQ_1_AN_SE_EQ_1 = 1.0,
       tsetup_posedge$D$CPN$CDN_EQ_1_AN_SE_EQ_0 = 1.0,
       thold_posedge$D$CPN$CDN_EQ_1_AN_SE_EQ_0 = 1.0,
       tsetup_posedge$SE$CPN$CDN_EQ_1 = 1.0,
       thold_posedge$SE$CPN$CDN_EQ_1 = 1.0,
       tsetup_posedge$SI$CPN$CDN_EQ_1_AN_SE_EQ_1 = 1.0,
       thold_posedge$SI$CPN$CDN_EQ_1_AN_SE_EQ_1 = 1.0,
       trec$CDN$CPN$D_EQ_0_AN_SE_EQ_1_AN_SI_EQ_1 = 1.0,
       trem$CDN$CPN$D_EQ_0_AN_SE_EQ_1_AN_SI_EQ_1 = 1.0;

     // path delays
     (negedge CPN *> (QN -: SE?SI:D)) = (tphlh$CPN$QN, tphhl$CPN$QN);
     (negedge CPN *> (Q +: SE?SI:D)) = (tphlh$CPN$Q, tphhl$CPN$Q);
     (negedge CDN *> (QN +: 1'b1)) = (tphlh$CDN$QN, 0);
     (negedge CDN *> (Q -: 1'b1)) = (0, tphhl$CDN$Q);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_SE_EQ_0 == 1'b1, negedge D, tsetup_negedge$D$CPN$CDN_EQ_1_AN_SE_EQ_0, thold_negedge$D$CPN$CDN_EQ_1_AN_SE_EQ_0, NOTIFIER);
     $setuphold(negedge CPN &&& CDN == 1'b1, negedge SE, tsetup_negedge$SE$CPN$CDN_EQ_1, thold_negedge$SE$CPN$CDN_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_SE_EQ_1 == 1'b1, negedge SI, tsetup_negedge$SI$CPN$CDN_EQ_1_AN_SE_EQ_1, thold_negedge$SI$CPN$CDN_EQ_1_AN_SE_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_SE_EQ_0 == 1'b1, posedge D, tsetup_posedge$D$CPN$CDN_EQ_1_AN_SE_EQ_0, thold_posedge$D$CPN$CDN_EQ_1_AN_SE_EQ_0, NOTIFIER);
     $setuphold(negedge CPN &&& CDN == 1'b1, posedge SE, tsetup_posedge$SE$CPN$CDN_EQ_1, thold_posedge$SE$CPN$CDN_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_SE_EQ_1 == 1'b1, posedge SI, tsetup_posedge$SI$CPN$CDN_EQ_1_AN_SE_EQ_1, thold_posedge$SI$CPN$CDN_EQ_1_AN_SE_EQ_1, NOTIFIER);
     $recrem(posedge CDN, negedge CPN &&& D_EQ_0_AN_SE_EQ_1_AN_SI_EQ_1 == 1'b1, trec$CDN$CPN$D_EQ_0_AN_SE_EQ_1_AN_SI_EQ_1, trem$CDN$CPN$D_EQ_0_AN_SE_EQ_1_AN_SI_EQ_1, NOTIFIER);
     $width(negedge CDN &&& D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$CDN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(posedge CPN &&& CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwh$CPN$CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(negedge CPN &&& CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$CPN$CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_SDF06D4 (Q, QN, CDN, CPN, D, SE, SI);
input  CDN ;
input  CPN ;
input  D ;
input  SE ;
input  SI ;
output Q ;
output QN ;
reg NOTIFIER ;

   udp_mux2 (I0_D, D, SI, SE);
   not (I0_CLOCK, CPN);
   not (I0_CLEAR, CDN);
   udp_dff (N_S_XM31_G, I0_D, I0_CLOCK, I0_CLEAR, 1'B0, NOTIFIER);
   not (N_NET0130_XM28_D, N_S_XM31_G);
   buf (Q, N_S_XM31_G);
   not (QN, N_S_XM31_G);
   and (CDN_EQ_1_AN_SE_EQ_1, CDN, SE);
   not (I10_out, SE);
   and (CDN_EQ_1_AN_SE_EQ_0, CDN, I10_out);
   not (I12_out, D);
   and (D_EQ_0_AN_SE_EQ_1_AN_SI_EQ_1, I12_out, SE, SI);
   not (I15_out, D);
   not (I16_out, SE);
   not (I18_out, SI);
   and (D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, I15_out, I16_out, I18_out);
   not (I20_out, D);
   not (I22_out, SE);
   not (I24_out, SI);
   and (CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, CDN, I20_out, I22_out, I24_out);

   specify
     // delay parameters
     specparam
       tphhl$CDN$Q = 1.0,
       tphlh$CDN$QN = 1.0,
       tphlh$CPN$Q = 1.0,
       tphhl$CPN$Q = 1.0,
       tphlh$CPN$QN = 1.0,
       tphhl$CPN$QN = 1.0,
       tminpwl$CDN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwh$CPN$CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwl$CPN$CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tsetup_negedge$D$CPN$CDN_EQ_1_AN_SE_EQ_0 = 1.0,
       thold_negedge$D$CPN$CDN_EQ_1_AN_SE_EQ_0 = 1.0,
       tsetup_negedge$SE$CPN$CDN_EQ_1 = 1.0,
       thold_negedge$SE$CPN$CDN_EQ_1 = 1.0,
       tsetup_negedge$SI$CPN$CDN_EQ_1_AN_SE_EQ_1 = 1.0,
       thold_negedge$SI$CPN$CDN_EQ_1_AN_SE_EQ_1 = 1.0,
       tsetup_posedge$D$CPN$CDN_EQ_1_AN_SE_EQ_0 = 1.0,
       thold_posedge$D$CPN$CDN_EQ_1_AN_SE_EQ_0 = 1.0,
       tsetup_posedge$SE$CPN$CDN_EQ_1 = 1.0,
       thold_posedge$SE$CPN$CDN_EQ_1 = 1.0,
       tsetup_posedge$SI$CPN$CDN_EQ_1_AN_SE_EQ_1 = 1.0,
       thold_posedge$SI$CPN$CDN_EQ_1_AN_SE_EQ_1 = 1.0,
       trec$CDN$CPN$D_EQ_0_AN_SE_EQ_1_AN_SI_EQ_1 = 1.0,
       trem$CDN$CPN$D_EQ_0_AN_SE_EQ_1_AN_SI_EQ_1 = 1.0;

     // path delays
     (negedge CPN *> (QN -: SE?SI:D)) = (tphlh$CPN$QN, tphhl$CPN$QN);
     (negedge CPN *> (Q +: SE?SI:D)) = (tphlh$CPN$Q, tphhl$CPN$Q);
     (negedge CDN *> (QN +: 1'b1)) = (tphlh$CDN$QN, 0);
     (negedge CDN *> (Q -: 1'b1)) = (0, tphhl$CDN$Q);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_SE_EQ_0 == 1'b1, negedge D, tsetup_negedge$D$CPN$CDN_EQ_1_AN_SE_EQ_0, thold_negedge$D$CPN$CDN_EQ_1_AN_SE_EQ_0, NOTIFIER);
     $setuphold(negedge CPN &&& CDN == 1'b1, negedge SE, tsetup_negedge$SE$CPN$CDN_EQ_1, thold_negedge$SE$CPN$CDN_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_SE_EQ_1 == 1'b1, negedge SI, tsetup_negedge$SI$CPN$CDN_EQ_1_AN_SE_EQ_1, thold_negedge$SI$CPN$CDN_EQ_1_AN_SE_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_SE_EQ_0 == 1'b1, posedge D, tsetup_posedge$D$CPN$CDN_EQ_1_AN_SE_EQ_0, thold_posedge$D$CPN$CDN_EQ_1_AN_SE_EQ_0, NOTIFIER);
     $setuphold(negedge CPN &&& CDN == 1'b1, posedge SE, tsetup_posedge$SE$CPN$CDN_EQ_1, thold_posedge$SE$CPN$CDN_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_SE_EQ_1 == 1'b1, posedge SI, tsetup_posedge$SI$CPN$CDN_EQ_1_AN_SE_EQ_1, thold_posedge$SI$CPN$CDN_EQ_1_AN_SE_EQ_1, NOTIFIER);
     $recrem(posedge CDN, negedge CPN &&& D_EQ_0_AN_SE_EQ_1_AN_SI_EQ_1 == 1'b1, trec$CDN$CPN$D_EQ_0_AN_SE_EQ_1_AN_SI_EQ_1, trem$CDN$CPN$D_EQ_0_AN_SE_EQ_1_AN_SI_EQ_1, NOTIFIER);
     $width(negedge CDN &&& D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$CDN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(posedge CPN &&& CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwh$CPN$CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(negedge CPN &&& CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$CPN$CDN_EQ_1_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_SDF07D1 (Q, QN, CPN, D, SDN, SE, SI);
input  CPN ;
input  D ;
input  SDN ;
input  SE ;
input  SI ;
output Q ;
output QN ;
reg NOTIFIER ;

   udp_mux2 (I0_D, D, SI, SE);
   not (I0_CLOCK, CPN);
   not (I0_SET, SDN);
   udp_dff (N_S_XM29_G, I0_D, I0_CLOCK, 1'B0, I0_SET, NOTIFIER);
   not (N_NET0130_XM26_D, N_S_XM29_G);
   buf (Q, N_S_XM29_G);
   not (QN, N_S_XM29_G);
   and (SDN_EQ_1_AN_SE_EQ_1, SDN, SE);
   not (I10_out, D);
   not (I11_out, SE);
   not (I13_out, SI);
   and (D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, I10_out, I11_out, I13_out);
   not (I15_out, SE);
   and (SDN_EQ_1_AN_SE_EQ_0, SDN, I15_out);
   not (I17_out, D);
   not (I19_out, SE);
   not (I21_out, SI);
   and (D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, I17_out, SDN, I19_out, I21_out);

   specify
     // delay parameters
     specparam
       tphlh$CPN$Q = 1.0,
       tphhl$CPN$Q = 1.0,
       tphlh$CPN$QN = 1.0,
       tphhl$CPN$QN = 1.0,
       tphlh$SDN$Q = 1.0,
       tphhl$SDN$QN = 1.0,
       tminpwh$CPN$D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwl$CPN$D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwl$SDN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tsetup_negedge$D$CPN$SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       thold_negedge$D$CPN$SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       tsetup_negedge$SE$CPN$SDN_EQ_1 = 1.0,
       thold_negedge$SE$CPN$SDN_EQ_1 = 1.0,
       tsetup_negedge$SI$CPN$SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       thold_negedge$SI$CPN$SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       tsetup_posedge$D$CPN$SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       thold_posedge$D$CPN$SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       tsetup_posedge$SE$CPN$SDN_EQ_1 = 1.0,
       thold_posedge$SE$CPN$SDN_EQ_1 = 1.0,
       tsetup_posedge$SI$CPN$SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       thold_posedge$SI$CPN$SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       trec$SDN$CPN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       trem$SDN$CPN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0;

     // path delays
     (negedge CPN *> (QN -: SE?SI:D)) = (tphlh$CPN$QN, tphhl$CPN$QN);
     (negedge CPN *> (Q +: SE?SI:D)) = (tphlh$CPN$Q, tphhl$CPN$Q);
     (negedge SDN *> (QN -: 1'b1)) = (0, tphhl$SDN$QN);
     (negedge SDN *> (Q +: 1'b1)) = (tphlh$SDN$Q, 0);
     $setuphold(negedge CPN &&& SDN_EQ_1_AN_SE_EQ_0 == 1'b1, negedge D, tsetup_negedge$D$CPN$SDN_EQ_1_AN_SE_EQ_0, thold_negedge$D$CPN$SDN_EQ_1_AN_SE_EQ_0, NOTIFIER);
     $setuphold(negedge CPN &&& SDN == 1'b1, negedge SE, tsetup_negedge$SE$CPN$SDN_EQ_1, thold_negedge$SE$CPN$SDN_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& SDN_EQ_1_AN_SE_EQ_1 == 1'b1, negedge SI, tsetup_negedge$SI$CPN$SDN_EQ_1_AN_SE_EQ_1, thold_negedge$SI$CPN$SDN_EQ_1_AN_SE_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& SDN_EQ_1_AN_SE_EQ_0 == 1'b1, posedge D, tsetup_posedge$D$CPN$SDN_EQ_1_AN_SE_EQ_0, thold_posedge$D$CPN$SDN_EQ_1_AN_SE_EQ_0, NOTIFIER);
     $setuphold(negedge CPN &&& SDN == 1'b1, posedge SE, tsetup_posedge$SE$CPN$SDN_EQ_1, thold_posedge$SE$CPN$SDN_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& SDN_EQ_1_AN_SE_EQ_1 == 1'b1, posedge SI, tsetup_posedge$SI$CPN$SDN_EQ_1_AN_SE_EQ_1, thold_posedge$SI$CPN$SDN_EQ_1_AN_SE_EQ_1, NOTIFIER);
     $recrem(posedge SDN, negedge CPN &&& D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, trec$SDN$CPN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, trem$SDN$CPN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, NOTIFIER);
     $width(posedge CPN &&& D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwh$CPN$D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(negedge CPN &&& D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$CPN$D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(negedge SDN &&& D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$SDN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_SDF07D2 (Q, QN, CPN, D, SDN, SE, SI);
input  CPN ;
input  D ;
input  SDN ;
input  SE ;
input  SI ;
output Q ;
output QN ;
reg NOTIFIER ;

   udp_mux2 (I0_D, D, SI, SE);
   not (I0_CLOCK, CPN);
   not (I0_SET, SDN);
   udp_dff (N_S_XM29_G, I0_D, I0_CLOCK, 1'B0, I0_SET, NOTIFIER);
   not (N_NET0130_XM26_D, N_S_XM29_G);
   buf (Q, N_S_XM29_G);
   not (QN, N_S_XM29_G);
   and (SDN_EQ_1_AN_SE_EQ_1, SDN, SE);
   not (I10_out, D);
   not (I11_out, SE);
   not (I13_out, SI);
   and (D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, I10_out, I11_out, I13_out);
   not (I15_out, SE);
   and (SDN_EQ_1_AN_SE_EQ_0, SDN, I15_out);
   not (I17_out, D);
   not (I19_out, SE);
   not (I21_out, SI);
   and (D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, I17_out, SDN, I19_out, I21_out);

   specify
     // delay parameters
     specparam
       tphlh$CPN$Q = 1.0,
       tphhl$CPN$Q = 1.0,
       tphlh$CPN$QN = 1.0,
       tphhl$CPN$QN = 1.0,
       tphlh$SDN$Q = 1.0,
       tphhl$SDN$QN = 1.0,
       tminpwh$CPN$D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwl$CPN$D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwl$SDN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tsetup_negedge$D$CPN$SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       thold_negedge$D$CPN$SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       tsetup_negedge$SE$CPN$SDN_EQ_1 = 1.0,
       thold_negedge$SE$CPN$SDN_EQ_1 = 1.0,
       tsetup_negedge$SI$CPN$SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       thold_negedge$SI$CPN$SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       tsetup_posedge$D$CPN$SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       thold_posedge$D$CPN$SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       tsetup_posedge$SE$CPN$SDN_EQ_1 = 1.0,
       thold_posedge$SE$CPN$SDN_EQ_1 = 1.0,
       tsetup_posedge$SI$CPN$SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       thold_posedge$SI$CPN$SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       trec$SDN$CPN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       trem$SDN$CPN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0;

     // path delays
     (negedge CPN *> (QN -: SE?SI:D)) = (tphlh$CPN$QN, tphhl$CPN$QN);
     (negedge CPN *> (Q +: SE?SI:D)) = (tphlh$CPN$Q, tphhl$CPN$Q);
     (negedge SDN *> (QN -: 1'b1)) = (0, tphhl$SDN$QN);
     (negedge SDN *> (Q +: 1'b1)) = (tphlh$SDN$Q, 0);
     $setuphold(negedge CPN &&& SDN_EQ_1_AN_SE_EQ_0 == 1'b1, negedge D, tsetup_negedge$D$CPN$SDN_EQ_1_AN_SE_EQ_0, thold_negedge$D$CPN$SDN_EQ_1_AN_SE_EQ_0, NOTIFIER);
     $setuphold(negedge CPN &&& SDN == 1'b1, negedge SE, tsetup_negedge$SE$CPN$SDN_EQ_1, thold_negedge$SE$CPN$SDN_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& SDN_EQ_1_AN_SE_EQ_1 == 1'b1, negedge SI, tsetup_negedge$SI$CPN$SDN_EQ_1_AN_SE_EQ_1, thold_negedge$SI$CPN$SDN_EQ_1_AN_SE_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& SDN_EQ_1_AN_SE_EQ_0 == 1'b1, posedge D, tsetup_posedge$D$CPN$SDN_EQ_1_AN_SE_EQ_0, thold_posedge$D$CPN$SDN_EQ_1_AN_SE_EQ_0, NOTIFIER);
     $setuphold(negedge CPN &&& SDN == 1'b1, posedge SE, tsetup_posedge$SE$CPN$SDN_EQ_1, thold_posedge$SE$CPN$SDN_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& SDN_EQ_1_AN_SE_EQ_1 == 1'b1, posedge SI, tsetup_posedge$SI$CPN$SDN_EQ_1_AN_SE_EQ_1, thold_posedge$SI$CPN$SDN_EQ_1_AN_SE_EQ_1, NOTIFIER);
     $recrem(posedge SDN, negedge CPN &&& D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, trec$SDN$CPN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, trem$SDN$CPN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, NOTIFIER);
     $width(posedge CPN &&& D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwh$CPN$D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(negedge CPN &&& D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$CPN$D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(negedge SDN &&& D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$SDN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_SDF07D4 (Q, QN, CPN, D, SDN, SE, SI);
input  CPN ;
input  D ;
input  SDN ;
input  SE ;
input  SI ;
output Q ;
output QN ;
reg NOTIFIER ;

   udp_mux2 (I0_D, D, SI, SE);
   not (I0_CLOCK, CPN);
   not (I0_SET, SDN);
   udp_dff (N_S_XM29_G, I0_D, I0_CLOCK, 1'B0, I0_SET, NOTIFIER);
   not (N_NET0130_XM26_D, N_S_XM29_G);
   buf (Q, N_S_XM29_G);
   not (QN, N_S_XM29_G);
   and (SDN_EQ_1_AN_SE_EQ_1, SDN, SE);
   not (I10_out, D);
   not (I11_out, SE);
   not (I13_out, SI);
   and (D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, I10_out, I11_out, I13_out);
   not (I15_out, SE);
   and (SDN_EQ_1_AN_SE_EQ_0, SDN, I15_out);
   not (I17_out, D);
   not (I19_out, SE);
   not (I21_out, SI);
   and (D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, I17_out, SDN, I19_out, I21_out);

   specify
     // delay parameters
     specparam
       tphlh$CPN$Q = 1.0,
       tphhl$CPN$Q = 1.0,
       tphlh$CPN$QN = 1.0,
       tphhl$CPN$QN = 1.0,
       tphlh$SDN$Q = 1.0,
       tphhl$SDN$QN = 1.0,
       tminpwh$CPN$D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwl$CPN$D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwl$SDN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tsetup_negedge$D$CPN$SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       thold_negedge$D$CPN$SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       tsetup_negedge$SE$CPN$SDN_EQ_1 = 1.0,
       thold_negedge$SE$CPN$SDN_EQ_1 = 1.0,
       tsetup_negedge$SI$CPN$SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       thold_negedge$SI$CPN$SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       tsetup_posedge$D$CPN$SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       thold_posedge$D$CPN$SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       tsetup_posedge$SE$CPN$SDN_EQ_1 = 1.0,
       thold_posedge$SE$CPN$SDN_EQ_1 = 1.0,
       tsetup_posedge$SI$CPN$SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       thold_posedge$SI$CPN$SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       trec$SDN$CPN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       trem$SDN$CPN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0;

     // path delays
     (negedge CPN *> (QN -: SE?SI:D)) = (tphlh$CPN$QN, tphhl$CPN$QN);
     (negedge CPN *> (Q +: SE?SI:D)) = (tphlh$CPN$Q, tphhl$CPN$Q);
     (negedge SDN *> (QN -: 1'b1)) = (0, tphhl$SDN$QN);
     (negedge SDN *> (Q +: 1'b1)) = (tphlh$SDN$Q, 0);
     $setuphold(negedge CPN &&& SDN_EQ_1_AN_SE_EQ_0 == 1'b1, negedge D, tsetup_negedge$D$CPN$SDN_EQ_1_AN_SE_EQ_0, thold_negedge$D$CPN$SDN_EQ_1_AN_SE_EQ_0, NOTIFIER);
     $setuphold(negedge CPN &&& SDN == 1'b1, negedge SE, tsetup_negedge$SE$CPN$SDN_EQ_1, thold_negedge$SE$CPN$SDN_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& SDN_EQ_1_AN_SE_EQ_1 == 1'b1, negedge SI, tsetup_negedge$SI$CPN$SDN_EQ_1_AN_SE_EQ_1, thold_negedge$SI$CPN$SDN_EQ_1_AN_SE_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& SDN_EQ_1_AN_SE_EQ_0 == 1'b1, posedge D, tsetup_posedge$D$CPN$SDN_EQ_1_AN_SE_EQ_0, thold_posedge$D$CPN$SDN_EQ_1_AN_SE_EQ_0, NOTIFIER);
     $setuphold(negedge CPN &&& SDN == 1'b1, posedge SE, tsetup_posedge$SE$CPN$SDN_EQ_1, thold_posedge$SE$CPN$SDN_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& SDN_EQ_1_AN_SE_EQ_1 == 1'b1, posedge SI, tsetup_posedge$SI$CPN$SDN_EQ_1_AN_SE_EQ_1, thold_posedge$SI$CPN$SDN_EQ_1_AN_SE_EQ_1, NOTIFIER);
     $recrem(posedge SDN, negedge CPN &&& D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, trec$SDN$CPN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, trem$SDN$CPN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, NOTIFIER);
     $width(posedge CPN &&& D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwh$CPN$D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(negedge CPN &&& D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$CPN$D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(negedge SDN &&& D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$SDN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_SDF08D1 (Q, QN, CDN, CPN, D, SDN, SE, SI);
input  CDN ;
input  CPN ;
input  D ;
input  SDN ;
input  SE ;
input  SI ;
output Q ;
output QN ;
reg NOTIFIER ;

   udp_mux2 (I0_D, D, SI, SE);
   not (I0_CLOCK, CPN);
   not (I0_CLEAR, CDN);
   not (I0_SET, SDN);
   udp_dff (N_S_XM33_G, I0_D, I0_CLOCK, I0_CLEAR, I0_SET, NOTIFIER);
   not (N_NET0130_XM30_D, N_S_XM33_G);
   not (Q, N_NET0130_XM30_D);
   buf (QN, N_NET0130_XM30_D);
   and (CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1, CDN, SDN, SE);
   and (CDN_EQ_1_AN_SDN_EQ_1, CDN, SDN);
   not (I14_out, SE);
   and (CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0, CDN, SDN, I14_out);
   not (I16_out, D);
   not (I17_out, SE);
   not (I19_out, SI);
   and (D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, I16_out, I17_out, I19_out);
   not (I21_out, D);
   not (I23_out, SE);
   not (I25_out, SI);
   and (D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, I21_out, SDN, I23_out, I25_out);
   not (I27_out, D);
   not (I30_out, SE);
   not (I32_out, SI);
   and (CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, CDN, I27_out, SDN, I30_out, I32_out);
   not (I34_out, CDN);
   not (I35_out, D);
   not (I37_out, SE);
   not (I39_out, SI);
   and (CDN_EQ_0_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, I34_out, I35_out, I37_out, I39_out);

   specify
     // delay parameters
     specparam
       tphhl$CDN$Q = 1.0,
       tphlh$CDN$QN = 1.0,
       tphlh$CPN$Q = 1.0,
       tphhl$CPN$Q = 1.0,
       tphlh$CPN$QN = 1.0,
       tphhl$CPN$QN = 1.0,
       tplhl$SDN$Q = 1.0,
       tphlh$SDN$Q = 1.0,
       tpllh$SDN$QN = 1.0,
       tphhl$SDN$QN = 1.0,
       tminpwl$CDN$D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwh$CPN$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwl$CPN$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwl$SDN$CDN_EQ_0_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tsetup_negedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       thold_negedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       tsetup_negedge$SE$CPN$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       thold_negedge$SE$CPN$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       tsetup_negedge$SI$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       thold_negedge$SI$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       tsetup_posedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       thold_posedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       tsetup_posedge$SE$CPN$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       thold_posedge$SE$CPN$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       tsetup_posedge$SI$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       thold_posedge$SI$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       trec$CDN$CPN$SDN_EQ_1 = 1.0,
       trem$CDN$CPN$SDN_EQ_1 = 1.0,
       trec$CDN$SDN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       trec$SDN$CPN$CDN_EQ_1 = 1.0,
       trem$SDN$CPN$CDN_EQ_1 = 1.0;

     // path delays
     (negedge CPN *> (QN -: SE?SI:D)) = (tphlh$CPN$QN, tphhl$CPN$QN);
     (negedge CPN *> (Q +: SE?SI:D)) = (tphlh$CPN$Q, tphhl$CPN$Q);
     (negedge SDN *> (QN -: 1'b1)) = (tpllh$SDN$QN, tphhl$SDN$QN);
     (negedge SDN *> (Q +: 1'b1)) = (tphlh$SDN$Q, tplhl$SDN$Q);
     (negedge CDN *> (QN +: 1'b1)) = (tphlh$CDN$QN, 0);
     (negedge CDN *> (Q -: 1'b1)) = (0, tphhl$CDN$Q);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0 == 1'b1, negedge D, tsetup_negedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0, thold_negedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0, NOTIFIER);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_SDN_EQ_1 == 1'b1, negedge SE, tsetup_negedge$SE$CPN$CDN_EQ_1_AN_SDN_EQ_1, thold_negedge$SE$CPN$CDN_EQ_1_AN_SDN_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1 == 1'b1, negedge SI, tsetup_negedge$SI$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1, thold_negedge$SI$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0 == 1'b1, posedge D, tsetup_posedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0, thold_posedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0, NOTIFIER);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_SDN_EQ_1 == 1'b1, posedge SE, tsetup_posedge$SE$CPN$CDN_EQ_1_AN_SDN_EQ_1, thold_posedge$SE$CPN$CDN_EQ_1_AN_SDN_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1 == 1'b1, posedge SI, tsetup_posedge$SI$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1, thold_posedge$SI$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1, NOTIFIER);
     $recrem(posedge CDN, negedge CPN &&& SDN == 1'b1, trec$CDN$CPN$SDN_EQ_1, trem$CDN$CPN$SDN_EQ_1, NOTIFIER);
     $recovery(posedge CDN, posedge SDN &&& D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, trec$CDN$SDN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, NOTIFIER);
     $recrem(posedge SDN, negedge CPN &&& CDN == 1'b1, trec$SDN$CPN$CDN_EQ_1, trem$SDN$CPN$CDN_EQ_1, NOTIFIER);
     $width(negedge CDN &&& D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$CDN$D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(posedge CPN &&& CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwh$CPN$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(negedge CPN &&& CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$CPN$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(negedge SDN &&& CDN_EQ_0_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$SDN$CDN_EQ_0_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_SDF08D2 (Q, QN, CDN, CPN, D, SDN, SE, SI);
input  CDN ;
input  CPN ;
input  D ;
input  SDN ;
input  SE ;
input  SI ;
output Q ;
output QN ;
reg NOTIFIER ;

   udp_mux2 (I0_D, D, SI, SE);
   not (I0_CLOCK, CPN);
   not (I0_CLEAR, CDN);
   not (I0_SET, SDN);
   udp_dff (N_S_XM33_G, I0_D, I0_CLOCK, I0_CLEAR, I0_SET, NOTIFIER);
   not (N_NET0130_XM30_D, N_S_XM33_G);
   not (Q, N_NET0130_XM30_D);
   buf (QN, N_NET0130_XM30_D);
   and (CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1, CDN, SDN, SE);
   and (CDN_EQ_1_AN_SDN_EQ_1, CDN, SDN);
   not (I14_out, SE);
   and (CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0, CDN, SDN, I14_out);
   not (I16_out, D);
   not (I17_out, SE);
   not (I19_out, SI);
   and (D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, I16_out, I17_out, I19_out);
   not (I21_out, D);
   not (I23_out, SE);
   not (I25_out, SI);
   and (D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, I21_out, SDN, I23_out, I25_out);
   not (I27_out, D);
   not (I30_out, SE);
   not (I32_out, SI);
   and (CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, CDN, I27_out, SDN, I30_out, I32_out);
   not (I34_out, CDN);
   not (I35_out, D);
   not (I37_out, SE);
   not (I39_out, SI);
   and (CDN_EQ_0_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, I34_out, I35_out, I37_out, I39_out);

   specify
     // delay parameters
     specparam
       tphhl$CDN$Q = 1.0,
       tphlh$CDN$QN = 1.0,
       tphlh$CPN$Q = 1.0,
       tphhl$CPN$Q = 1.0,
       tphlh$CPN$QN = 1.0,
       tphhl$CPN$QN = 1.0,
       tplhl$SDN$Q = 1.0,
       tphlh$SDN$Q = 1.0,
       tpllh$SDN$QN = 1.0,
       tphhl$SDN$QN = 1.0,
       tminpwl$CDN$D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwh$CPN$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwl$CPN$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwl$SDN$CDN_EQ_0_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tsetup_negedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       thold_negedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       tsetup_negedge$SE$CPN$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       thold_negedge$SE$CPN$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       tsetup_negedge$SI$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       thold_negedge$SI$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       tsetup_posedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       thold_posedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       tsetup_posedge$SE$CPN$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       thold_posedge$SE$CPN$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       tsetup_posedge$SI$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       thold_posedge$SI$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       trec$CDN$CPN$SDN_EQ_1 = 1.0,
       trem$CDN$CPN$SDN_EQ_1 = 1.0,
       trec$CDN$SDN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       trec$SDN$CPN$CDN_EQ_1 = 1.0,
       trem$SDN$CPN$CDN_EQ_1 = 1.0;

     // path delays
     (negedge CPN *> (QN -: SE?SI:D)) = (tphlh$CPN$QN, tphhl$CPN$QN);
     (negedge CPN *> (Q +: SE?SI:D)) = (tphlh$CPN$Q, tphhl$CPN$Q);
     (negedge SDN *> (QN -: 1'b1)) = (tpllh$SDN$QN, tphhl$SDN$QN);
     (negedge SDN *> (Q +: 1'b1)) = (tphlh$SDN$Q, tplhl$SDN$Q);
     (negedge CDN *> (QN +: 1'b1)) = (tphlh$CDN$QN, 0);
     (negedge CDN *> (Q -: 1'b1)) = (0, tphhl$CDN$Q);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0 == 1'b1, negedge D, tsetup_negedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0, thold_negedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0, NOTIFIER);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_SDN_EQ_1 == 1'b1, negedge SE, tsetup_negedge$SE$CPN$CDN_EQ_1_AN_SDN_EQ_1, thold_negedge$SE$CPN$CDN_EQ_1_AN_SDN_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1 == 1'b1, negedge SI, tsetup_negedge$SI$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1, thold_negedge$SI$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0 == 1'b1, posedge D, tsetup_posedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0, thold_posedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0, NOTIFIER);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_SDN_EQ_1 == 1'b1, posedge SE, tsetup_posedge$SE$CPN$CDN_EQ_1_AN_SDN_EQ_1, thold_posedge$SE$CPN$CDN_EQ_1_AN_SDN_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1 == 1'b1, posedge SI, tsetup_posedge$SI$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1, thold_posedge$SI$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1, NOTIFIER);
     $recrem(posedge CDN, negedge CPN &&& SDN == 1'b1, trec$CDN$CPN$SDN_EQ_1, trem$CDN$CPN$SDN_EQ_1, NOTIFIER);
     $recovery(posedge CDN, posedge SDN &&& D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, trec$CDN$SDN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, NOTIFIER);
     $recrem(posedge SDN, negedge CPN &&& CDN == 1'b1, trec$SDN$CPN$CDN_EQ_1, trem$SDN$CPN$CDN_EQ_1, NOTIFIER);
     $width(negedge CDN &&& D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$CDN$D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(posedge CPN &&& CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwh$CPN$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(negedge CPN &&& CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$CPN$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(negedge SDN &&& CDN_EQ_0_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$SDN$CDN_EQ_0_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_SDF08D4 (Q, QN, CDN, CPN, D, SDN, SE, SI);
input  CDN ;
input  CPN ;
input  D ;
input  SDN ;
input  SE ;
input  SI ;
output Q ;
output QN ;
reg NOTIFIER ;

   udp_mux2 (I0_D, D, SI, SE);
   not (I0_CLOCK, CPN);
   not (I0_CLEAR, CDN);
   not (I0_SET, SDN);
   udp_dff (N_S_XM33_G, I0_D, I0_CLOCK, I0_CLEAR, I0_SET, NOTIFIER);
   not (N_NET0130_XM30_D, N_S_XM33_G);
   not (Q, N_NET0130_XM30_D);
   buf (QN, N_NET0130_XM30_D);
   and (CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1, CDN, SDN, SE);
   and (CDN_EQ_1_AN_SDN_EQ_1, CDN, SDN);
   not (I14_out, SE);
   and (CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0, CDN, SDN, I14_out);
   not (I16_out, D);
   not (I17_out, SE);
   not (I19_out, SI);
   and (D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, I16_out, I17_out, I19_out);
   not (I21_out, D);
   not (I23_out, SE);
   not (I25_out, SI);
   and (D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, I21_out, SDN, I23_out, I25_out);
   not (I27_out, D);
   not (I30_out, SE);
   not (I32_out, SI);
   and (CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, CDN, I27_out, SDN, I30_out, I32_out);
   not (I34_out, CDN);
   not (I35_out, D);
   not (I37_out, SE);
   not (I39_out, SI);
   and (CDN_EQ_0_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, I34_out, I35_out, I37_out, I39_out);

   specify
     // delay parameters
     specparam
       tphhl$CDN$Q = 1.0,
       tphlh$CDN$QN = 1.0,
       tphlh$CPN$Q = 1.0,
       tphhl$CPN$Q = 1.0,
       tphlh$CPN$QN = 1.0,
       tphhl$CPN$QN = 1.0,
       tplhl$SDN$Q = 1.0,
       tphlh$SDN$Q = 1.0,
       tpllh$SDN$QN = 1.0,
       tphhl$SDN$QN = 1.0,
       tminpwl$CDN$D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwh$CPN$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwl$CPN$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tminpwl$SDN$CDN_EQ_0_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       tsetup_negedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       thold_negedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       tsetup_negedge$SE$CPN$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       thold_negedge$SE$CPN$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       tsetup_negedge$SI$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       thold_negedge$SI$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       tsetup_posedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       thold_posedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0 = 1.0,
       tsetup_posedge$SE$CPN$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       thold_posedge$SE$CPN$CDN_EQ_1_AN_SDN_EQ_1 = 1.0,
       tsetup_posedge$SI$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       thold_posedge$SI$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1 = 1.0,
       trec$CDN$CPN$SDN_EQ_1 = 1.0,
       trem$CDN$CPN$SDN_EQ_1 = 1.0,
       trec$CDN$SDN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 = 1.0,
       trec$SDN$CPN$CDN_EQ_1 = 1.0,
       trem$SDN$CPN$CDN_EQ_1 = 1.0;

     // path delays
     (negedge CPN *> (QN -: SE?SI:D)) = (tphlh$CPN$QN, tphhl$CPN$QN);
     (negedge CPN *> (Q +: SE?SI:D)) = (tphlh$CPN$Q, tphhl$CPN$Q);
     (negedge SDN *> (QN -: 1'b1)) = (tpllh$SDN$QN, tphhl$SDN$QN);
     (negedge SDN *> (Q +: 1'b1)) = (tphlh$SDN$Q, tplhl$SDN$Q);
     (negedge CDN *> (QN +: 1'b1)) = (tphlh$CDN$QN, 0);
     (negedge CDN *> (Q -: 1'b1)) = (0, tphhl$CDN$Q);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0 == 1'b1, negedge D, tsetup_negedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0, thold_negedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0, NOTIFIER);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_SDN_EQ_1 == 1'b1, negedge SE, tsetup_negedge$SE$CPN$CDN_EQ_1_AN_SDN_EQ_1, thold_negedge$SE$CPN$CDN_EQ_1_AN_SDN_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1 == 1'b1, negedge SI, tsetup_negedge$SI$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1, thold_negedge$SI$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0 == 1'b1, posedge D, tsetup_posedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0, thold_posedge$D$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_0, NOTIFIER);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_SDN_EQ_1 == 1'b1, posedge SE, tsetup_posedge$SE$CPN$CDN_EQ_1_AN_SDN_EQ_1, thold_posedge$SE$CPN$CDN_EQ_1_AN_SDN_EQ_1, NOTIFIER);
     $setuphold(negedge CPN &&& CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1 == 1'b1, posedge SI, tsetup_posedge$SI$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1, thold_posedge$SI$CPN$CDN_EQ_1_AN_SDN_EQ_1_AN_SE_EQ_1, NOTIFIER);
     $recrem(posedge CDN, negedge CPN &&& SDN == 1'b1, trec$CDN$CPN$SDN_EQ_1, trem$CDN$CPN$SDN_EQ_1, NOTIFIER);
     $recovery(posedge CDN, posedge SDN &&& D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, trec$CDN$SDN$D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, NOTIFIER);
     $recrem(posedge SDN, negedge CPN &&& CDN == 1'b1, trec$SDN$CPN$CDN_EQ_1, trem$SDN$CPN$CDN_EQ_1, NOTIFIER);
     $width(negedge CDN &&& D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$CDN$D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(posedge CPN &&& CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwh$CPN$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(negedge CPN &&& CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$CPN$CDN_EQ_1_AN_D_EQ_0_AN_SDN_EQ_1_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);
     $width(negedge SDN &&& CDN_EQ_0_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0 == 1'b1, tminpwl$SDN$CDN_EQ_0_AN_D_EQ_0_AN_SE_EQ_0_AN_SI_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_TL01D1 (ECK, CK, E);
input  CK ;
input  E ;
output ECK ;
reg NOTIFIER ;
reg ReSeT;

`ifdef  RSTn_lib
	 initial begin
		ReSeT = 0 ;
		#3 ReSeT = 1 ;
		#111 ReSeT = 0 ;
	end
  `else initial  ReSeT = 0;
`endif

   not (I0_ENABLE, CK);
   udp_tlat (N_NM_XM9_G, E, I0_ENABLE, ReSeT /*1'B0*/, 1'B0, NOTIFIER);
   not (N_M_XM6_D, N_NM_XM9_G);
   and (ECK, CK, N_NM_XM9_G);

   specify
     // delay parameters
     specparam
       tpllh$CK$ECK = 1.0,
       tphhl$CK$ECK = 1.0,
       tminpwl$CK$E_EQ_0 = 1.0,
       tsetup_negedge$E$CK = 1.0,
       thold_negedge$E$CK = 1.0,
       tsetup_posedge$E$CK = 1.0,
       thold_posedge$E$CK = 1.0;

     // path delays
     (posedge CK *> (ECK +: 1'b1)) = (tpllh$CK$ECK, 0);
     (negedge CK *> (ECK -: 1'b1)) = (0, tphhl$CK$ECK);
     $setuphold(posedge CK, negedge E, tsetup_negedge$E$CK, thold_negedge$E$CK, NOTIFIER);
     $setuphold(posedge CK, posedge E, tsetup_posedge$E$CK, thold_posedge$E$CK, NOTIFIER);
     $width(negedge CK &&& E == 1'b0, tminpwl$CK$E_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_TL01D2 (ECK, CK, E);
input  CK ;
input  E ;
output ECK ;
reg NOTIFIER ;
reg ReSeT;

`ifdef  RSTn_lib
	 initial begin
		ReSeT = 0 ;
		#3 ReSeT = 1 ;
		#111 ReSeT = 0 ;
	end
  `else initial  ReSeT = 0;
`endif

   not (I0_ENABLE, CK);
   udp_tlat (N_NM_XM9_G, E, I0_ENABLE,  ReSeT /*1'B0*/, 1'B0, NOTIFIER);
   not (N_M_XM6_D, N_NM_XM9_G);
   and (ECK, CK, N_NM_XM9_G);

   specify
     // delay parameters
     specparam
       tpllh$CK$ECK = 1.0,
       tphhl$CK$ECK = 1.0,
       tminpwl$CK$E_EQ_0 = 1.0,
       tsetup_negedge$E$CK = 1.0,
       thold_negedge$E$CK = 1.0,
       tsetup_posedge$E$CK = 1.0,
       thold_posedge$E$CK = 1.0;

     // path delays
     (posedge CK *> (ECK +: 1'b1)) = (tpllh$CK$ECK, 0);
     (negedge CK *> (ECK -: 1'b1)) = (0, tphhl$CK$ECK);
     $setuphold(posedge CK, negedge E, tsetup_negedge$E$CK, thold_negedge$E$CK, NOTIFIER);
     $setuphold(posedge CK, posedge E, tsetup_posedge$E$CK, thold_posedge$E$CK, NOTIFIER);
     $width(negedge CK &&& E == 1'b0, tminpwl$CK$E_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_TL01D4 (ECK, CK, E);
input  CK ;
input  E ;
output ECK ;
reg NOTIFIER ;
reg ReSeT;

`ifdef  RSTn_lib
	 initial begin
		ReSeT = 0 ;
		#3 ReSeT = 1 ;
		#111 ReSeT = 0 ;
	end
  `else initial  ReSeT = 0;
`endif

   not (I0_ENABLE, CK);
   udp_tlat (N_NM_XM9_G, E, I0_ENABLE,  ReSeT /*1'B0*/, 1'B0, NOTIFIER);
   not (N_M_XM6_D, N_NM_XM9_G);
   and (ECK, CK, N_NM_XM9_G);

   specify
     // delay parameters
     specparam
       tpllh$CK$ECK = 1.0,
       tphhl$CK$ECK = 1.0,
       tminpwl$CK$E_EQ_0 = 1.0,
       tsetup_negedge$E$CK = 1.0,
       thold_negedge$E$CK = 1.0,
       tsetup_posedge$E$CK = 1.0,
       thold_posedge$E$CK = 1.0;

     // path delays
     (posedge CK *> (ECK +: 1'b1)) = (tpllh$CK$ECK, 0);
     (negedge CK *> (ECK -: 1'b1)) = (0, tphhl$CK$ECK);
     $setuphold(posedge CK, negedge E, tsetup_negedge$E$CK, thold_negedge$E$CK, NOTIFIER);
     $setuphold(posedge CK, posedge E, tsetup_posedge$E$CK, thold_posedge$E$CK, NOTIFIER);
     $width(negedge CK &&& E == 1'b0, tminpwl$CK$E_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_TL01D6 (ECK, CK, E);
input  CK ;
input  E ;
output ECK ;
reg NOTIFIER ;
// _ILJA_
reg ReSeT;

`ifdef  RSTn_lib
	 initial begin
		ReSeT = 0 ;
		#3 ReSeT = 1 ;
		#111 ReSeT = 0 ;
	end
  `else initial  ReSeT = 0;
`endif

   not (I0_ENABLE, CK);
   udp_tlat (N_NM_XM15_G, E, I0_ENABLE, ReSeT/*1'B0*/, 1'B0, NOTIFIER);
   not (N_M_XM6_D, N_NM_XM15_G);
   and (ECK, CK, N_NM_XM15_G);

   specify
     // delay parameters
     specparam
       tpllh$CK$ECK = 1.0,
       tphhl$CK$ECK = 1.0,
       tminpwl$CK$E_EQ_0 = 1.0,
       tsetup_negedge$E$CK = 1.0,
       thold_negedge$E$CK = 1.0,
       tsetup_posedge$E$CK = 1.0,
       thold_posedge$E$CK = 1.0;

     // path delays
     (posedge CK *> (ECK +: 1'b1)) = (tpllh$CK$ECK, 0);
     (negedge CK *> (ECK -: 1'b1)) = (0, tphhl$CK$ECK);
     $setuphold(posedge CK, negedge E, tsetup_negedge$E$CK, thold_negedge$E$CK, NOTIFIER);
     $setuphold(posedge CK, posedge E, tsetup_posedge$E$CK, thold_posedge$E$CK, NOTIFIER);
     $width(negedge CK &&& E == 1'b0, tminpwl$CK$E_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_TL01D8 (ECK, CK, E);
input  CK ;
input  E ;
output ECK ;
reg NOTIFIER ;
reg ReSeT;


`ifdef  RSTn_lib
	 initial begin
		ReSeT = 0 ;
		#3 ReSeT = 1 ;
		#111 ReSeT = 0 ;
	end
  `else initial  ReSeT = 0;
`endif

   not (I0_ENABLE, CK);
  udp_tlat (N_NM_XM15_G, E, I0_ENABLE,  ReSeT /*1'B0*/, 1'B0, NOTIFIER);
   not (N_M_XM6_D, N_NM_XM15_G);
   and (ECK, CK, N_NM_XM15_G);

   specify
     // delay parameters
     specparam
       tpllh$CK$ECK = 1.0,
       tphhl$CK$ECK = 1.0,
       tminpwl$CK$E_EQ_0 = 1.0,
       tsetup_negedge$E$CK = 1.0,
       thold_negedge$E$CK = 1.0,
       tsetup_posedge$E$CK = 1.0,
       thold_posedge$E$CK = 1.0;

     // path delays
     (posedge CK *> (ECK +: 1'b1)) = (tpllh$CK$ECK, 0);
     (negedge CK *> (ECK -: 1'b1)) = (0, tphhl$CK$ECK);
     $setuphold(posedge CK, negedge E, tsetup_negedge$E$CK, thold_negedge$E$CK, NOTIFIER);
     $setuphold(posedge CK, posedge E, tsetup_posedge$E$CK, thold_posedge$E$CK, NOTIFIER);
     $width(negedge CK &&& E == 1'b0, tminpwl$CK$E_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_TL02D1 (ECKN, CKN, E);
input  CKN ;
input  E ;
output ECKN ;
reg NOTIFIER ;

   udp_tlat (N_NM_XM9_G, E, CKN, 1'B0, 1'B0, NOTIFIER);
   not (N_M_XM17_G, N_NM_XM9_G);
   or  (ECKN, CKN, N_M_XM17_G);

   specify
     // delay parameters
     specparam
       tpllh$CKN$ECKN = 1.0,
       tphhl$CKN$ECKN = 1.0,
       tminpwh$CKN$E_EQ_0 = 1.0,
       tsetup_negedge$E$CKN = 1.0,
       thold_negedge$E$CKN = 1.0,
       tsetup_posedge$E$CKN = 1.0,
       thold_posedge$E$CKN = 1.0;

     // path delays
     (posedge CKN *> (ECKN +: 1'b1)) = (tpllh$CKN$ECKN, 0);
     (negedge CKN *> (ECKN -: 1'b1)) = (0, tphhl$CKN$ECKN);
     $setuphold(negedge CKN, negedge E, tsetup_negedge$E$CKN, thold_negedge$E$CKN, NOTIFIER);
     $setuphold(negedge CKN, posedge E, tsetup_posedge$E$CKN, thold_posedge$E$CKN, NOTIFIER);
     $width(posedge CKN &&& E == 1'b0, tminpwh$CKN$E_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_TL02D2 (ECKN, CKN, E);
input  CKN ;
input  E ;
output ECKN ;
reg NOTIFIER ;

   udp_tlat (N_NM_XM9_G, E, CKN, 1'B0, 1'B0, NOTIFIER);
   not (N_M_XM17_G, N_NM_XM9_G);
   or  (ECKN, CKN, N_M_XM17_G);

   specify
     // delay parameters
     specparam
       tpllh$CKN$ECKN = 1.0,
       tphhl$CKN$ECKN = 1.0,
       tminpwh$CKN$E_EQ_0 = 1.0,
       tsetup_negedge$E$CKN = 1.0,
       thold_negedge$E$CKN = 1.0,
       tsetup_posedge$E$CKN = 1.0,
       thold_posedge$E$CKN = 1.0;

     // path delays
     (posedge CKN *> (ECKN +: 1'b1)) = (tpllh$CKN$ECKN, 0);
     (negedge CKN *> (ECKN -: 1'b1)) = (0, tphhl$CKN$ECKN);
     $setuphold(negedge CKN, negedge E, tsetup_negedge$E$CKN, thold_negedge$E$CKN, NOTIFIER);
     $setuphold(negedge CKN, posedge E, tsetup_posedge$E$CKN, thold_posedge$E$CKN, NOTIFIER);
     $width(posedge CKN &&& E == 1'b0, tminpwh$CKN$E_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_TL02D4 (ECKN, CKN, E);
input  CKN ;
input  E ;
output ECKN ;
reg NOTIFIER ;

   udp_tlat (N_NM_XM9_G, E, CKN, 1'B0, 1'B0, NOTIFIER);
   not (N_M_XM17_G, N_NM_XM9_G);
   or  (ECKN, CKN, N_M_XM17_G);

   specify
     // delay parameters
     specparam
       tpllh$CKN$ECKN = 1.0,
       tphhl$CKN$ECKN = 1.0,
       tminpwh$CKN$E_EQ_0 = 1.0,
       tsetup_negedge$E$CKN = 1.0,
       thold_negedge$E$CKN = 1.0,
       tsetup_posedge$E$CKN = 1.0,
       thold_posedge$E$CKN = 1.0;

     // path delays
     (posedge CKN *> (ECKN +: 1'b1)) = (tpllh$CKN$ECKN, 0);
     (negedge CKN *> (ECKN -: 1'b1)) = (0, tphhl$CKN$ECKN);
     $setuphold(negedge CKN, negedge E, tsetup_negedge$E$CKN, thold_negedge$E$CKN, NOTIFIER);
     $setuphold(negedge CKN, posedge E, tsetup_posedge$E$CKN, thold_posedge$E$CKN, NOTIFIER);
     $width(posedge CKN &&& E == 1'b0, tminpwh$CKN$E_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_TL03D1 (ECK, CK, E, SE);
input  CK ;
input  E ;
input  SE ;
output ECK ;
reg NOTIFIER ;

   or  (I0_D, E, SE);
   not (I0_ENABLE, CK);
   udp_tlat (N_NM_XM11_G, I0_D, I0_ENABLE, 1'B0, 1'B0, NOTIFIER);
   not (N_M_XM7_D, N_NM_XM11_G);
   and (ECK, CK, N_NM_XM11_G);
   not (I6_out, E);
   not (I7_out, SE);
   and (E_EQ_0_AN_SE_EQ_0, I6_out, I7_out);

   specify
     // delay parameters
     specparam
       tpllh$CK$ECK = 1.0,
       tphhl$CK$ECK = 1.0,
       tminpwl$CK$E_EQ_0_AN_SE_EQ_0 = 1.0,
       tsetup_negedge$E$CK$SE_EQ_0 = 1.0,
       thold_negedge$E$CK$SE_EQ_0 = 1.0,
       tsetup_negedge$SE$CK$E_EQ_0 = 1.0,
       thold_negedge$SE$CK$E_EQ_0 = 1.0,
       tsetup_posedge$E$CK$SE_EQ_0 = 1.0,
       thold_posedge$E$CK$SE_EQ_0 = 1.0,
       tsetup_posedge$SE$CK$E_EQ_0 = 1.0,
       thold_posedge$SE$CK$E_EQ_0 = 1.0;

     // path delays
     (posedge CK *> (ECK +: 1'b1)) = (tpllh$CK$ECK, 0);
     (negedge CK *> (ECK -: 1'b1)) = (0, tphhl$CK$ECK);
     $setuphold(posedge CK &&& SE == 1'b0, negedge E, tsetup_negedge$E$CK$SE_EQ_0, thold_negedge$E$CK$SE_EQ_0, NOTIFIER);
     $setuphold(posedge CK &&& E == 1'b0, negedge SE, tsetup_negedge$SE$CK$E_EQ_0, thold_negedge$SE$CK$E_EQ_0, NOTIFIER);
     $setuphold(posedge CK &&& SE == 1'b0, posedge E, tsetup_posedge$E$CK$SE_EQ_0, thold_posedge$E$CK$SE_EQ_0, NOTIFIER);
     $setuphold(posedge CK &&& E == 1'b0, posedge SE, tsetup_posedge$SE$CK$E_EQ_0, thold_posedge$SE$CK$E_EQ_0, NOTIFIER);
     $width(negedge CK &&& E_EQ_0_AN_SE_EQ_0 == 1'b1, tminpwl$CK$E_EQ_0_AN_SE_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_TL03D2 (ECK, CK, E, SE);
input  CK ;
input  E ;
input  SE ;
output ECK ;
reg NOTIFIER ;

   or  (I0_D, E, SE);
   not (I0_ENABLE, CK);
   udp_tlat (N_NM_XM11_G, I0_D, I0_ENABLE, 1'B0, 1'B0, NOTIFIER);
   not (N_M_XM7_D, N_NM_XM11_G);
   and (ECK, CK, N_NM_XM11_G);
   not (I6_out, E);
   not (I7_out, SE);
   and (E_EQ_0_AN_SE_EQ_0, I6_out, I7_out);

   specify
     // delay parameters
     specparam
       tpllh$CK$ECK = 1.0,
       tphhl$CK$ECK = 1.0,
       tminpwl$CK$E_EQ_0_AN_SE_EQ_0 = 1.0,
       tsetup_negedge$E$CK$SE_EQ_0 = 1.0,
       thold_negedge$E$CK$SE_EQ_0 = 1.0,
       tsetup_negedge$SE$CK$E_EQ_0 = 1.0,
       thold_negedge$SE$CK$E_EQ_0 = 1.0,
       tsetup_posedge$E$CK$SE_EQ_0 = 1.0,
       thold_posedge$E$CK$SE_EQ_0 = 1.0,
       tsetup_posedge$SE$CK$E_EQ_0 = 1.0,
       thold_posedge$SE$CK$E_EQ_0 = 1.0;

     // path delays
     (posedge CK *> (ECK +: 1'b1)) = (tpllh$CK$ECK, 0);
     (negedge CK *> (ECK -: 1'b1)) = (0, tphhl$CK$ECK);
     $setuphold(posedge CK &&& SE == 1'b0, negedge E, tsetup_negedge$E$CK$SE_EQ_0, thold_negedge$E$CK$SE_EQ_0, NOTIFIER);
     $setuphold(posedge CK &&& E == 1'b0, negedge SE, tsetup_negedge$SE$CK$E_EQ_0, thold_negedge$SE$CK$E_EQ_0, NOTIFIER);
     $setuphold(posedge CK &&& SE == 1'b0, posedge E, tsetup_posedge$E$CK$SE_EQ_0, thold_posedge$E$CK$SE_EQ_0, NOTIFIER);
     $setuphold(posedge CK &&& E == 1'b0, posedge SE, tsetup_posedge$SE$CK$E_EQ_0, thold_posedge$SE$CK$E_EQ_0, NOTIFIER);
     $width(negedge CK &&& E_EQ_0_AN_SE_EQ_0 == 1'b1, tminpwl$CK$E_EQ_0_AN_SE_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_TL03D4 (ECK, CK, E, SE);
input  CK ;
input  E ;
input  SE ;
output ECK ;
reg NOTIFIER ;

   or  (I0_D, E, SE);
   not (I0_ENABLE, CK);
   udp_tlat (N_NM_XM11_G, I0_D, I0_ENABLE, 1'B0, 1'B0, NOTIFIER);
   not (N_M_XM7_D, N_NM_XM11_G);
   and (ECK, CK, N_NM_XM11_G);
   not (I6_out, E);
   not (I7_out, SE);
   and (E_EQ_0_AN_SE_EQ_0, I6_out, I7_out);

   specify
     // delay parameters
     specparam
       tpllh$CK$ECK = 1.0,
       tphhl$CK$ECK = 1.0,
       tminpwl$CK$E_EQ_0_AN_SE_EQ_0 = 1.0,
       tsetup_negedge$E$CK$SE_EQ_0 = 1.0,
       thold_negedge$E$CK$SE_EQ_0 = 1.0,
       tsetup_negedge$SE$CK$E_EQ_0 = 1.0,
       thold_negedge$SE$CK$E_EQ_0 = 1.0,
       tsetup_posedge$E$CK$SE_EQ_0 = 1.0,
       thold_posedge$E$CK$SE_EQ_0 = 1.0,
       tsetup_posedge$SE$CK$E_EQ_0 = 1.0,
       thold_posedge$SE$CK$E_EQ_0 = 1.0;

     // path delays
     (posedge CK *> (ECK +: 1'b1)) = (tpllh$CK$ECK, 0);
     (negedge CK *> (ECK -: 1'b1)) = (0, tphhl$CK$ECK);
     $setuphold(posedge CK &&& SE == 1'b0, negedge E, tsetup_negedge$E$CK$SE_EQ_0, thold_negedge$E$CK$SE_EQ_0, NOTIFIER);
     $setuphold(posedge CK &&& E == 1'b0, negedge SE, tsetup_negedge$SE$CK$E_EQ_0, thold_negedge$SE$CK$E_EQ_0, NOTIFIER);
     $setuphold(posedge CK &&& SE == 1'b0, posedge E, tsetup_posedge$E$CK$SE_EQ_0, thold_posedge$E$CK$SE_EQ_0, NOTIFIER);
     $setuphold(posedge CK &&& E == 1'b0, posedge SE, tsetup_posedge$SE$CK$E_EQ_0, thold_posedge$SE$CK$E_EQ_0, NOTIFIER);
     $width(negedge CK &&& E_EQ_0_AN_SE_EQ_0 == 1'b1, tminpwl$CK$E_EQ_0_AN_SE_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_TL03D6 (ECK, CK, E, SE);
input  CK ;
input  E ;
input  SE ;
output ECK ;
reg NOTIFIER ;

   or  (I0_D, E, SE);
   not (I0_ENABLE, CK);
   udp_tlat (N_NM_XM11_G, I0_D, I0_ENABLE, 1'B0, 1'B0, NOTIFIER);
   not (N_M_XM7_D, N_NM_XM11_G);
   and (ECK, CK, N_NM_XM11_G);
   not (I6_out, E);
   not (I7_out, SE);
   and (E_EQ_0_AN_SE_EQ_0, I6_out, I7_out);

   specify
     // delay parameters
     specparam
       tpllh$CK$ECK = 1.0,
       tphhl$CK$ECK = 1.0,
       tminpwl$CK$E_EQ_0_AN_SE_EQ_0 = 1.0,
       tsetup_negedge$E$CK$SE_EQ_0 = 1.0,
       thold_negedge$E$CK$SE_EQ_0 = 1.0,
       tsetup_negedge$SE$CK$E_EQ_0 = 1.0,
       thold_negedge$SE$CK$E_EQ_0 = 1.0,
       tsetup_posedge$E$CK$SE_EQ_0 = 1.0,
       thold_posedge$E$CK$SE_EQ_0 = 1.0,
       tsetup_posedge$SE$CK$E_EQ_0 = 1.0,
       thold_posedge$SE$CK$E_EQ_0 = 1.0;

     // path delays
     (posedge CK *> (ECK +: 1'b1)) = (tpllh$CK$ECK, 0);
     (negedge CK *> (ECK -: 1'b1)) = (0, tphhl$CK$ECK);
     $setuphold(posedge CK &&& SE == 1'b0, negedge E, tsetup_negedge$E$CK$SE_EQ_0, thold_negedge$E$CK$SE_EQ_0, NOTIFIER);
     $setuphold(posedge CK &&& E == 1'b0, negedge SE, tsetup_negedge$SE$CK$E_EQ_0, thold_negedge$SE$CK$E_EQ_0, NOTIFIER);
     $setuphold(posedge CK &&& SE == 1'b0, posedge E, tsetup_posedge$E$CK$SE_EQ_0, thold_posedge$E$CK$SE_EQ_0, NOTIFIER);
     $setuphold(posedge CK &&& E == 1'b0, posedge SE, tsetup_posedge$SE$CK$E_EQ_0, thold_posedge$SE$CK$E_EQ_0, NOTIFIER);
     $width(negedge CK &&& E_EQ_0_AN_SE_EQ_0 == 1'b1, tminpwl$CK$E_EQ_0_AN_SE_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_TL03D8 (ECK, CK, E, SE);
input  CK ;
input  E ;
input  SE ;
output ECK ;
reg NOTIFIER ;

   or  (I0_D, E, SE);
   not (I0_ENABLE, CK);
   udp_tlat (N_NM_XM11_G, I0_D, I0_ENABLE, 1'B0, 1'B0, NOTIFIER);
   not (N_M_XM7_D, N_NM_XM11_G);
   and (ECK, CK, N_NM_XM11_G);
   not (I6_out, E);
   not (I7_out, SE);
   and (E_EQ_0_AN_SE_EQ_0, I6_out, I7_out);

   specify
     // delay parameters
     specparam
       tpllh$CK$ECK = 1.0,
       tphhl$CK$ECK = 1.0,
       tminpwl$CK$E_EQ_0_AN_SE_EQ_0 = 1.0,
       tsetup_negedge$E$CK$SE_EQ_0 = 1.0,
       thold_negedge$E$CK$SE_EQ_0 = 1.0,
       tsetup_negedge$SE$CK$E_EQ_0 = 1.0,
       thold_negedge$SE$CK$E_EQ_0 = 1.0,
       tsetup_posedge$E$CK$SE_EQ_0 = 1.0,
       thold_posedge$E$CK$SE_EQ_0 = 1.0,
       tsetup_posedge$SE$CK$E_EQ_0 = 1.0,
       thold_posedge$SE$CK$E_EQ_0 = 1.0;

     // path delays
     (posedge CK *> (ECK +: 1'b1)) = (tpllh$CK$ECK, 0);
     (negedge CK *> (ECK -: 1'b1)) = (0, tphhl$CK$ECK);
     $setuphold(posedge CK &&& SE == 1'b0, negedge E, tsetup_negedge$E$CK$SE_EQ_0, thold_negedge$E$CK$SE_EQ_0, NOTIFIER);
     $setuphold(posedge CK &&& E == 1'b0, negedge SE, tsetup_negedge$SE$CK$E_EQ_0, thold_negedge$SE$CK$E_EQ_0, NOTIFIER);
     $setuphold(posedge CK &&& SE == 1'b0, posedge E, tsetup_posedge$E$CK$SE_EQ_0, thold_posedge$E$CK$SE_EQ_0, NOTIFIER);
     $setuphold(posedge CK &&& E == 1'b0, posedge SE, tsetup_posedge$SE$CK$E_EQ_0, thold_posedge$SE$CK$E_EQ_0, NOTIFIER);
     $width(negedge CK &&& E_EQ_0_AN_SE_EQ_0 == 1'b1, tminpwl$CK$E_EQ_0_AN_SE_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_TL04D1 (ECKN, CKN, E, SE);
input  CKN ;
input  E ;
input  SE ;
output ECKN ;
reg NOTIFIER ;

   or  (I0_D, E, SE);
   udp_tlat (N_NM_XM11_G, I0_D, CKN, 1'B0, 1'B0, NOTIFIER);
   not (N_M_XM7_D, N_NM_XM11_G);
   or  (ECKN, CKN, N_M_XM7_D);
   not (I5_out, E);
   not (I6_out, SE);
   and (E_EQ_0_AN_SE_EQ_0, I5_out, I6_out);

   specify
     // delay parameters
     specparam
       tpllh$CKN$ECKN = 1.0,
       tphhl$CKN$ECKN = 1.0,
       tminpwh$CKN$E_EQ_0_AN_SE_EQ_0 = 1.0,
       tsetup_negedge$E$CKN$SE_EQ_0 = 1.0,
       thold_negedge$E$CKN$SE_EQ_0 = 1.0,
       tsetup_negedge$SE$CKN$E_EQ_0 = 1.0,
       thold_negedge$SE$CKN$E_EQ_0 = 1.0,
       tsetup_posedge$E$CKN$SE_EQ_0 = 1.0,
       thold_posedge$E$CKN$SE_EQ_0 = 1.0,
       tsetup_posedge$SE$CKN$E_EQ_0 = 1.0,
       thold_posedge$SE$CKN$E_EQ_0 = 1.0;

     // path delays
     (posedge CKN *> (ECKN +: 1'b1)) = (tpllh$CKN$ECKN, 0);
     (negedge CKN *> (ECKN -: 1'b1)) = (0, tphhl$CKN$ECKN);
     $setuphold(negedge CKN &&& SE == 1'b0, negedge E, tsetup_negedge$E$CKN$SE_EQ_0, thold_negedge$E$CKN$SE_EQ_0, NOTIFIER);
     $setuphold(negedge CKN &&& E == 1'b0, negedge SE, tsetup_negedge$SE$CKN$E_EQ_0, thold_negedge$SE$CKN$E_EQ_0, NOTIFIER);
     $setuphold(negedge CKN &&& SE == 1'b0, posedge E, tsetup_posedge$E$CKN$SE_EQ_0, thold_posedge$E$CKN$SE_EQ_0, NOTIFIER);
     $setuphold(negedge CKN &&& E == 1'b0, posedge SE, tsetup_posedge$SE$CKN$E_EQ_0, thold_posedge$SE$CKN$E_EQ_0, NOTIFIER);
     $width(posedge CKN &&& E_EQ_0_AN_SE_EQ_0 == 1'b1, tminpwh$CKN$E_EQ_0_AN_SE_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_TL04D2 (ECKN, CKN, E, SE);
input  CKN ;
input  E ;
input  SE ;
output ECKN ;
reg NOTIFIER ;

   or  (I0_D, E, SE);
   udp_tlat (N_NM_XM11_G, I0_D, CKN, 1'B0, 1'B0, NOTIFIER);
   not (N_M_XM7_D, N_NM_XM11_G);
   or  (ECKN, CKN, N_M_XM7_D);
   not (I5_out, E);
   not (I6_out, SE);
   and (E_EQ_0_AN_SE_EQ_0, I5_out, I6_out);

   specify
     // delay parameters
     specparam
       tpllh$CKN$ECKN = 1.0,
       tphhl$CKN$ECKN = 1.0,
       tminpwh$CKN$E_EQ_0_AN_SE_EQ_0 = 1.0,
       tsetup_negedge$E$CKN$SE_EQ_0 = 1.0,
       thold_negedge$E$CKN$SE_EQ_0 = 1.0,
       tsetup_negedge$SE$CKN$E_EQ_0 = 1.0,
       thold_negedge$SE$CKN$E_EQ_0 = 1.0,
       tsetup_posedge$E$CKN$SE_EQ_0 = 1.0,
       thold_posedge$E$CKN$SE_EQ_0 = 1.0,
       tsetup_posedge$SE$CKN$E_EQ_0 = 1.0,
       thold_posedge$SE$CKN$E_EQ_0 = 1.0;

     // path delays
     (posedge CKN *> (ECKN +: 1'b1)) = (tpllh$CKN$ECKN, 0);
     (negedge CKN *> (ECKN -: 1'b1)) = (0, tphhl$CKN$ECKN);
     $setuphold(negedge CKN &&& SE == 1'b0, negedge E, tsetup_negedge$E$CKN$SE_EQ_0, thold_negedge$E$CKN$SE_EQ_0, NOTIFIER);
     $setuphold(negedge CKN &&& E == 1'b0, negedge SE, tsetup_negedge$SE$CKN$E_EQ_0, thold_negedge$SE$CKN$E_EQ_0, NOTIFIER);
     $setuphold(negedge CKN &&& SE == 1'b0, posedge E, tsetup_posedge$E$CKN$SE_EQ_0, thold_posedge$E$CKN$SE_EQ_0, NOTIFIER);
     $setuphold(negedge CKN &&& E == 1'b0, posedge SE, tsetup_posedge$SE$CKN$E_EQ_0, thold_posedge$SE$CKN$E_EQ_0, NOTIFIER);
     $width(posedge CKN &&& E_EQ_0_AN_SE_EQ_0 == 1'b1, tminpwh$CKN$E_EQ_0_AN_SE_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_TL04D4 (ECKN, CKN, E, SE);
input  CKN ;
input  E ;
input  SE ;
output ECKN ;
reg NOTIFIER ;

   or  (I0_D, E, SE);
   udp_tlat (N_NM_XM11_G, I0_D, CKN, 1'B0, 1'B0, NOTIFIER);
   not (N_M_XM7_D, N_NM_XM11_G);
   or  (ECKN, CKN, N_M_XM7_D);
   not (I5_out, E);
   not (I6_out, SE);
   and (E_EQ_0_AN_SE_EQ_0, I5_out, I6_out);

   specify
     // delay parameters
     specparam
       tpllh$CKN$ECKN = 1.0,
       tphhl$CKN$ECKN = 1.0,
       tminpwh$CKN$E_EQ_0_AN_SE_EQ_0 = 1.0,
       tsetup_negedge$E$CKN$SE_EQ_0 = 1.0,
       thold_negedge$E$CKN$SE_EQ_0 = 1.0,
       tsetup_negedge$SE$CKN$E_EQ_0 = 1.0,
       thold_negedge$SE$CKN$E_EQ_0 = 1.0,
       tsetup_posedge$E$CKN$SE_EQ_0 = 1.0,
       thold_posedge$E$CKN$SE_EQ_0 = 1.0,
       tsetup_posedge$SE$CKN$E_EQ_0 = 1.0,
       thold_posedge$SE$CKN$E_EQ_0 = 1.0;

     // path delays
     (posedge CKN *> (ECKN +: 1'b1)) = (tpllh$CKN$ECKN, 0);
     (negedge CKN *> (ECKN -: 1'b1)) = (0, tphhl$CKN$ECKN);
     $setuphold(negedge CKN &&& SE == 1'b0, negedge E, tsetup_negedge$E$CKN$SE_EQ_0, thold_negedge$E$CKN$SE_EQ_0, NOTIFIER);
     $setuphold(negedge CKN &&& E == 1'b0, negedge SE, tsetup_negedge$SE$CKN$E_EQ_0, thold_negedge$SE$CKN$E_EQ_0, NOTIFIER);
     $setuphold(negedge CKN &&& SE == 1'b0, posedge E, tsetup_posedge$E$CKN$SE_EQ_0, thold_posedge$E$CKN$SE_EQ_0, NOTIFIER);
     $setuphold(negedge CKN &&& E == 1'b0, posedge SE, tsetup_posedge$SE$CKN$E_EQ_0, thold_posedge$SE$CKN$E_EQ_0, NOTIFIER);
     $width(posedge CKN &&& E_EQ_0_AN_SE_EQ_0 == 1'b1, tminpwh$CKN$E_EQ_0_AN_SE_EQ_0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_XN02D1 (ZN, A1, A2);
input  A1 ;
input  A2 ;
output ZN ;

   xor (I0_out, A1, A2);
   not (ZN, I0_out);

   specify
     // delay parameters
     specparam
       tpllh$A1$ZN = 1.0,
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tphhl$A1$ZN = 1.0,
       tpllh$A2$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tphhl$A2$ZN = 1.0;

     // path delays
     (posedge A2 *> (ZN +: A1)) = (tpllh$A2$ZN, tplhl$A2$ZN);
     (negedge A2 *> (ZN +: !A1)) = (tphlh$A2$ZN, tphhl$A2$ZN);
     (posedge A1 *> (ZN +: A2)) = (tpllh$A1$ZN, tplhl$A1$ZN);
     (negedge A1 *> (ZN +: !A2)) = (tphlh$A1$ZN, tphhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_XN02D2 (ZN, A1, A2);
input  A1 ;
input  A2 ;
output ZN ;

   xor (I0_out, A1, A2);
   not (ZN, I0_out);

   specify
     // delay parameters
     specparam
       tpllh$A1$ZN = 1.0,
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tphhl$A1$ZN = 1.0,
       tpllh$A2$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tphhl$A2$ZN = 1.0;

     // path delays
     (posedge A2 *> (ZN +: A1)) = (tpllh$A2$ZN, tplhl$A2$ZN);
     (negedge A2 *> (ZN +: !A1)) = (tphlh$A2$ZN, tphhl$A2$ZN);
     (posedge A1 *> (ZN +: A2)) = (tpllh$A1$ZN, tplhl$A1$ZN);
     (negedge A1 *> (ZN +: !A2)) = (tphlh$A1$ZN, tphhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_XN02D4 (ZN, A1, A2);
input  A1 ;
input  A2 ;
output ZN ;

   xor (I0_out, A1, A2);
   not (ZN, I0_out);

   specify
     // delay parameters
     specparam
       tpllh$A1$ZN = 1.0,
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tphhl$A1$ZN = 1.0,
       tpllh$A2$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tphhl$A2$ZN = 1.0;

     // path delays
     (posedge A2 *> (ZN +: A1)) = (tpllh$A2$ZN, tplhl$A2$ZN);
     (negedge A2 *> (ZN +: !A1)) = (tphlh$A2$ZN, tphhl$A2$ZN);
     (posedge A1 *> (ZN +: A2)) = (tpllh$A1$ZN, tplhl$A1$ZN);
     (negedge A1 *> (ZN +: !A2)) = (tphlh$A1$ZN, tphhl$A1$ZN);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_XN03D1 (ZN, A1, A2, A3);
input  A1 ;
input  A2 ;
input  A3 ;
output ZN ;

   xor (I0_out, A1, A2);
   xor (I1_out, I0_out, A3);
   not (ZN, I1_out);

   specify
     // delay parameters
    /* specparam
       tpllh$A1$ZN = 1.0,
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tphhl$A1$ZN = 1.0,
       tpllh$A2$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tphhl$A2$ZN = 1.0,
       tpllh$A3$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0,
       tphhl$A3$ZN = 1.0,
       tpllh$A1$ZN$A2_EQ_0_AN_A3_EQ_1 = 1.0,
       tphhl$A1$ZN$A2_EQ_0_AN_A3_EQ_1 = 1.0,
       tpllh$A1$ZN$A2_EQ_1_AN_A3_EQ_0 = 1.0,
       tphhl$A1$ZN$A2_EQ_1_AN_A3_EQ_0 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0 = 1.0,
       tpllh$A2$ZN$A1_EQ_0_AN_A3_EQ_1 = 1.0,
       tphhl$A2$ZN$A1_EQ_0_AN_A3_EQ_1 = 1.0,
       tpllh$A2$ZN$A1_EQ_1_AN_A3_EQ_0 = 1.0,
       tphhl$A2$ZN$A1_EQ_1_AN_A3_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0 = 1.0,
       tpllh$A3$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0,
       tphhl$A3$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0,
       tpllh$A3$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tphhl$A3$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1 = 1.0,
       tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1 = 1.0,
       tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0 = 1.0,
       tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1, tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0)
       (A3 *> ZN) = (tpllh$A3$ZN$A1_EQ_1_AN_A2_EQ_0, tphhl$A3$ZN$A1_EQ_1_AN_A2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1)
       (A3 *> ZN) = (tpllh$A3$ZN$A1_EQ_0_AN_A2_EQ_1, tphhl$A3$ZN$A1_EQ_0_AN_A2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0, tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0);
     ifnone
       (A3 *> ZN) = (tpllh$A3$ZN,tplhl$A3$ZN);

     if (A1 == 1'b1 && A3 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1, tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1);
     if (A1 == 1'b1 && A3 == 1'b0)
       (A2 *> ZN) = (tpllh$A2$ZN$A1_EQ_1_AN_A3_EQ_0, tphhl$A2$ZN$A1_EQ_1_AN_A3_EQ_0);
     if (A1 == 1'b0 && A3 == 1'b1)
       (A2 *> ZN) = (tpllh$A2$ZN$A1_EQ_0_AN_A3_EQ_1, tphhl$A2$ZN$A1_EQ_0_AN_A3_EQ_1);
     if (A1 == 1'b0 && A3 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0, tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0);
     ifnone
       (A2 *> ZN) = (tpllh$A2$ZN,tplhl$A2$ZN);

     if (A2 == 1'b1 && A3 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1, tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1);
     if (A2 == 1'b1 && A3 == 1'b0)
       (A1 *> ZN) = (tpllh$A1$ZN$A2_EQ_1_AN_A3_EQ_0, tphhl$A1$ZN$A2_EQ_1_AN_A3_EQ_0);
     if (A2 == 1'b0 && A3 == 1'b1)
       (A1 *> ZN) = (tpllh$A1$ZN$A2_EQ_0_AN_A3_EQ_1, tphhl$A1$ZN$A2_EQ_0_AN_A3_EQ_1);
     if (A2 == 1'b0 && A3 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0, tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0);
     ifnone
       (A1 *> ZN) = (tpllh$A1$ZN,tplhl$A1$ZN);*/

 // path delays
      (posedge A1 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge A1 => (ZN -: ZN)) = (1.0, 1.0);
      if (A2 == 1'b0 && A3 == 1'b1) (A1 +=> ZN) = (1.0, 1.0);
      if (A2 == 1'b1 && A3 == 1'b0) (A1 +=> ZN) = (1.0, 1.0);
      if (A2 == 1'b1 && A3 == 1'b1) (A1 -=> ZN) = (1.0, 1.0);
      if (A2 == 1'b0 && A3 == 1'b0) (A1 -=> ZN) = (1.0, 1.0);


      (posedge A2 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge A2 => (ZN -: ZN)) = (1.0, 1.0);
      if (A1 == 1'b0 && A3 == 1'b1) (A2 +=> ZN) = (1.0, 1.0);
      if (A1 == 1'b1 && A3 == 1'b0) (A2 +=> ZN) = (1.0, 1.0);
      if (A1 == 1'b1 && A3 == 1'b1) (A2 -=> ZN) = (1.0, 1.0);
      if (A1 == 1'b0 && A3 == 1'b0) (A2 -=> ZN) = (1.0, 1.0);


      (posedge A3 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge A3 => (ZN -: ZN)) = (1.0, 1.0);
      if (A1 == 1'b1 && A2 == 1'b0) (A3 +=> ZN) = (1.0, 1.0);
      if (A1 == 1'b0 && A2 == 1'b1) (A3 +=> ZN) = (1.0, 1.0);
      if (A1 == 1'b1 && A2 == 1'b1) (A3 -=> ZN) = (1.0, 1.0);
      if (A1 == 1'b0 && A2 == 1'b0) (A3 -=> ZN) = (1.0, 1.0);



   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_XN03D2 (ZN, A1, A2, A3);
input  A1 ;
input  A2 ;
input  A3 ;
output ZN ;

   xor (I0_out, A1, A2);
   xor (I1_out, I0_out, A3);
   not (ZN, I1_out);

   specify
     // delay parameters
 /*    specparam
       tpllh$A1$ZN = 1.0,
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tphhl$A1$ZN = 1.0,
       tpllh$A2$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tphhl$A2$ZN = 1.0,
       tpllh$A3$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0,
       tphhl$A3$ZN = 1.0,
       tpllh$A1$ZN$A2_EQ_0_AN_A3_EQ_1 = 1.0,
       tphhl$A1$ZN$A2_EQ_0_AN_A3_EQ_1 = 1.0,
       tpllh$A1$ZN$A2_EQ_1_AN_A3_EQ_0 = 1.0,
       tphhl$A1$ZN$A2_EQ_1_AN_A3_EQ_0 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0 = 1.0,
       tpllh$A2$ZN$A1_EQ_0_AN_A3_EQ_1 = 1.0,
       tphhl$A2$ZN$A1_EQ_0_AN_A3_EQ_1 = 1.0,
       tpllh$A2$ZN$A1_EQ_1_AN_A3_EQ_0 = 1.0,
       tphhl$A2$ZN$A1_EQ_1_AN_A3_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0 = 1.0,
       tpllh$A3$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0,
       tphhl$A3$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0,
       tpllh$A3$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tphhl$A3$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1 = 1.0,
       tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1 = 1.0,
       tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0 = 1.0,
       tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1, tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0)
       (A3 *> ZN) = (tpllh$A3$ZN$A1_EQ_1_AN_A2_EQ_0, tphhl$A3$ZN$A1_EQ_1_AN_A2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1)
       (A3 *> ZN) = (tpllh$A3$ZN$A1_EQ_0_AN_A2_EQ_1, tphhl$A3$ZN$A1_EQ_0_AN_A2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0, tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0);
     ifnone
       (A3 *> ZN) = (tpllh$A3$ZN,tplhl$A3$ZN);

     if (A1 == 1'b1 && A3 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1, tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1);
     if (A1 == 1'b1 && A3 == 1'b0)
       (A2 *> ZN) = (tpllh$A2$ZN$A1_EQ_1_AN_A3_EQ_0, tphhl$A2$ZN$A1_EQ_1_AN_A3_EQ_0);
     if (A1 == 1'b0 && A3 == 1'b1)
       (A2 *> ZN) = (tpllh$A2$ZN$A1_EQ_0_AN_A3_EQ_1, tphhl$A2$ZN$A1_EQ_0_AN_A3_EQ_1);
     if (A1 == 1'b0 && A3 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0, tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0);
     ifnone
       (A2 *> ZN) = (tpllh$A2$ZN,tplhl$A2$ZN);

     if (A2 == 1'b1 && A3 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1, tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1);
     if (A2 == 1'b1 && A3 == 1'b0)
       (A1 *> ZN) = (tpllh$A1$ZN$A2_EQ_1_AN_A3_EQ_0, tphhl$A1$ZN$A2_EQ_1_AN_A3_EQ_0);
     if (A2 == 1'b0 && A3 == 1'b1)
       (A1 *> ZN) = (tpllh$A1$ZN$A2_EQ_0_AN_A3_EQ_1, tphhl$A1$ZN$A2_EQ_0_AN_A3_EQ_1);
     if (A2 == 1'b0 && A3 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0, tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0);
     ifnone
       (A1 *> ZN) = (tpllh$A1$ZN,tplhl$A1$ZN);*/
      (posedge A1 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge A1 => (ZN -: ZN)) = (1.0, 1.0);
      if (A2 == 1'b0 && A3 == 1'b1) (A1 +=> ZN) = (1.0, 1.0);
      if (A2 == 1'b1 && A3 == 1'b0) (A1 +=> ZN) = (1.0, 1.0);
      if (A2 == 1'b1 && A3 == 1'b1) (A1 -=> ZN) = (1.0, 1.0);
      if (A2 == 1'b0 && A3 == 1'b0) (A1 -=> ZN) = (1.0, 1.0);


      (posedge A2 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge A2 => (ZN -: ZN)) = (1.0, 1.0);
      if (A1 == 1'b0 && A3 == 1'b1) (A2 +=> ZN) = (1.0, 1.0);
      if (A1 == 1'b1 && A3 == 1'b0) (A2 +=> ZN) = (1.0, 1.0);
      if (A1 == 1'b1 && A3 == 1'b1) (A2 -=> ZN) = (1.0, 1.0);
      if (A1 == 1'b0 && A3 == 1'b0) (A2 -=> ZN) = (1.0, 1.0);


      (posedge A3 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge A3 => (ZN -: ZN)) = (1.0, 1.0);
      if (A1 == 1'b1 && A2 == 1'b0) (A3 +=> ZN) = (1.0, 1.0);
      if (A1 == 1'b0 && A2 == 1'b1) (A3 +=> ZN) = (1.0, 1.0);
      if (A1 == 1'b1 && A2 == 1'b1) (A3 -=> ZN) = (1.0, 1.0);
      if (A1 == 1'b0 && A2 == 1'b0) (A3 -=> ZN) = (1.0, 1.0);




   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_XN03D4 (ZN, A1, A2, A3);
input  A1 ;
input  A2 ;
input  A3 ;
output ZN ;

   xor (I0_out, A1, A2);
   xor (I1_out, I0_out, A3);
   not (ZN, I1_out);

   specify
     // delay parameters
 /*    specparam
       tpllh$A1$ZN = 1.0,
       tplhl$A1$ZN = 1.0,
       tphlh$A1$ZN = 1.0,
       tphhl$A1$ZN = 1.0,
       tpllh$A2$ZN = 1.0,
       tplhl$A2$ZN = 1.0,
       tphlh$A2$ZN = 1.0,
       tphhl$A2$ZN = 1.0,
       tpllh$A3$ZN = 1.0,
       tplhl$A3$ZN = 1.0,
       tphlh$A3$ZN = 1.0,
       tphhl$A3$ZN = 1.0,
       tpllh$A1$ZN$A2_EQ_0_AN_A3_EQ_1 = 1.0,
       tphhl$A1$ZN$A2_EQ_0_AN_A3_EQ_1 = 1.0,
       tpllh$A1$ZN$A2_EQ_1_AN_A3_EQ_0 = 1.0,
       tphhl$A1$ZN$A2_EQ_1_AN_A3_EQ_0 = 1.0,
       tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1 = 1.0,
       tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1 = 1.0,
       tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0 = 1.0,
       tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0 = 1.0,
       tpllh$A2$ZN$A1_EQ_0_AN_A3_EQ_1 = 1.0,
       tphhl$A2$ZN$A1_EQ_0_AN_A3_EQ_1 = 1.0,
       tpllh$A2$ZN$A1_EQ_1_AN_A3_EQ_0 = 1.0,
       tphhl$A2$ZN$A1_EQ_1_AN_A3_EQ_0 = 1.0,
       tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1 = 1.0,
       tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1 = 1.0,
       tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0 = 1.0,
       tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0 = 1.0,
       tpllh$A3$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0,
       tphhl$A3$ZN$A1_EQ_1_AN_A2_EQ_0 = 1.0,
       tpllh$A3$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tphhl$A3$ZN$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1 = 1.0,
       tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1 = 1.0,
       tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0 = 1.0,
       tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_1_AN_A2_EQ_1, tplhl$A3$ZN$A1_EQ_1_AN_A2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0)
       (A3 *> ZN) = (tpllh$A3$ZN$A1_EQ_1_AN_A2_EQ_0, tphhl$A3$ZN$A1_EQ_1_AN_A2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1)
       (A3 *> ZN) = (tpllh$A3$ZN$A1_EQ_0_AN_A2_EQ_1, tphhl$A3$ZN$A1_EQ_0_AN_A2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0)
       (A3 *> ZN) = (tphlh$A3$ZN$A1_EQ_0_AN_A2_EQ_0, tplhl$A3$ZN$A1_EQ_0_AN_A2_EQ_0);
     ifnone
       (A3 *> ZN) = (tpllh$A3$ZN,tplhl$A3$ZN);

     if (A1 == 1'b1 && A3 == 1'b1)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_1_AN_A3_EQ_1, tplhl$A2$ZN$A1_EQ_1_AN_A3_EQ_1);
     if (A1 == 1'b1 && A3 == 1'b0)
       (A2 *> ZN) = (tpllh$A2$ZN$A1_EQ_1_AN_A3_EQ_0, tphhl$A2$ZN$A1_EQ_1_AN_A3_EQ_0);
     if (A1 == 1'b0 && A3 == 1'b1)
       (A2 *> ZN) = (tpllh$A2$ZN$A1_EQ_0_AN_A3_EQ_1, tphhl$A2$ZN$A1_EQ_0_AN_A3_EQ_1);
     if (A1 == 1'b0 && A3 == 1'b0)
       (A2 *> ZN) = (tphlh$A2$ZN$A1_EQ_0_AN_A3_EQ_0, tplhl$A2$ZN$A1_EQ_0_AN_A3_EQ_0);
     ifnone
       (A2 *> ZN) = (tpllh$A2$ZN,tplhl$A2$ZN);

     if (A2 == 1'b1 && A3 == 1'b1)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_1_AN_A3_EQ_1, tplhl$A1$ZN$A2_EQ_1_AN_A3_EQ_1);
     if (A2 == 1'b1 && A3 == 1'b0)
       (A1 *> ZN) = (tpllh$A1$ZN$A2_EQ_1_AN_A3_EQ_0, tphhl$A1$ZN$A2_EQ_1_AN_A3_EQ_0);
     if (A2 == 1'b0 && A3 == 1'b1)
       (A1 *> ZN) = (tpllh$A1$ZN$A2_EQ_0_AN_A3_EQ_1, tphhl$A1$ZN$A2_EQ_0_AN_A3_EQ_1);
     if (A2 == 1'b0 && A3 == 1'b0)
       (A1 *> ZN) = (tphlh$A1$ZN$A2_EQ_0_AN_A3_EQ_0, tplhl$A1$ZN$A2_EQ_0_AN_A3_EQ_0);
     ifnone
       (A1 *> ZN) = (tpllh$A1$ZN,tplhl$A1$ZN);*/


     // path delays
      (posedge A1 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge A1 => (ZN -: ZN)) = (1.0, 1.0);
      if (A2 == 1'b0 && A3 == 1'b1) (A1 +=> ZN) = (1.0, 1.0);
      if (A2 == 1'b1 && A3 == 1'b0) (A1 +=> ZN) = (1.0, 1.0);
      if (A2 == 1'b1 && A3 == 1'b1) (A1 -=> ZN) = (1.0, 1.0);
      if (A2 == 1'b0 && A3 == 1'b0) (A1 -=> ZN) = (1.0, 1.0);


      (posedge A2 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge A2 => (ZN -: ZN)) = (1.0, 1.0);
      if (A1 == 1'b0 && A3 == 1'b1) (A2 +=> ZN) = (1.0, 1.0);
      if (A1 == 1'b1 && A3 == 1'b0) (A2 +=> ZN) = (1.0, 1.0);
      if (A1 == 1'b1 && A3 == 1'b1) (A2 -=> ZN) = (1.0, 1.0);
      if (A1 == 1'b0 && A3 == 1'b0) (A2 -=> ZN) = (1.0, 1.0);


      (posedge A3 => (ZN +: ZN)) = (1.0, 1.0);
      (negedge A3 => (ZN -: ZN)) = (1.0, 1.0);
      if (A1 == 1'b1 && A2 == 1'b0) (A3 +=> ZN) = (1.0, 1.0);
      if (A1 == 1'b0 && A2 == 1'b1) (A3 +=> ZN) = (1.0, 1.0);
      if (A1 == 1'b1 && A2 == 1'b1) (A3 -=> ZN) = (1.0, 1.0);
      if (A1 == 1'b0 && A2 == 1'b0) (A3 -=> ZN) = (1.0, 1.0);



   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_XO02D1 (Z, A1, A2);
input  A1 ;
input  A2 ;
output Z ;

   xor (Z, A1, A2);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tplhl$A1$Z = 1.0,
       tphlh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tplhl$A2$Z = 1.0,
       tphlh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0;

     // path delays
     (posedge A2 *> (Z +: !A1)) = (tpllh$A2$Z, tplhl$A2$Z);
     (negedge A2 *> (Z +: A1)) = (tphlh$A2$Z, tphhl$A2$Z);
     (posedge A1 *> (Z +: !A2)) = (tpllh$A1$Z, tplhl$A1$Z);
     (negedge A1 *> (Z +: A2)) = (tphlh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_XO02D2 (Z, A1, A2);
input  A1 ;
input  A2 ;
output Z ;

   xor (Z, A1, A2);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tplhl$A1$Z = 1.0,
       tphlh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tplhl$A2$Z = 1.0,
       tphlh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0;

     // path delays
     (posedge A2 *> (Z +: !A1)) = (tpllh$A2$Z, tplhl$A2$Z);
     (negedge A2 *> (Z +: A1)) = (tphlh$A2$Z, tphhl$A2$Z);
     (posedge A1 *> (Z +: !A2)) = (tpllh$A1$Z, tplhl$A1$Z);
     (negedge A1 *> (Z +: A2)) = (tphlh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_XO02D4 (Z, A1, A2);
input  A1 ;
input  A2 ;
output Z ;

   xor (Z, A1, A2);

   specify
     // delay parameters
     specparam
       tpllh$A1$Z = 1.0,
       tplhl$A1$Z = 1.0,
       tphlh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tplhl$A2$Z = 1.0,
       tphlh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0;

     // path delays
     (posedge A2 *> (Z +: !A1)) = (tpllh$A2$Z, tplhl$A2$Z);
     (negedge A2 *> (Z +: A1)) = (tphlh$A2$Z, tphhl$A2$Z);
     (posedge A1 *> (Z +: !A2)) = (tpllh$A1$Z, tplhl$A1$Z);
     (negedge A1 *> (Z +: A2)) = (tphlh$A1$Z, tphhl$A1$Z);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_XO03D1 (Z, A1, A2, A3);
input  A1 ;
input  A2 ;
input  A3 ;
output Z ;

   xor (I0_out, A1, A2);
   xor (Z, I0_out, A3);

   specify
     // delay parameters
   /*  specparam
       tpllh$A1$Z = 1.0,
       tplhl$A1$Z = 1.0,
       tphlh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tplhl$A2$Z = 1.0,
       tphlh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$A3$Z = 1.0,
       tplhl$A3$Z = 1.0,
       tphlh$A3$Z = 1.0,
       tphhl$A3$Z = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_A3_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_A3_EQ_1 = 1.0,
       tpllh$A1$Z$A2_EQ_0_AN_A3_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_0_AN_A3_EQ_0 = 1.0,
       tplhl$A1$Z$A2_EQ_0_AN_A3_EQ_1 = 1.0,
       tphlh$A1$Z$A2_EQ_0_AN_A3_EQ_1 = 1.0,
       tplhl$A1$Z$A2_EQ_1_AN_A3_EQ_0 = 1.0,
       tphlh$A1$Z$A2_EQ_1_AN_A3_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_A3_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_A3_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_0_AN_A3_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_0_AN_A3_EQ_0 = 1.0,
       tplhl$A2$Z$A1_EQ_0_AN_A3_EQ_1 = 1.0,
       tphlh$A2$Z$A1_EQ_0_AN_A3_EQ_1 = 1.0,
       tplhl$A2$Z$A1_EQ_1_AN_A3_EQ_0 = 1.0,
       tphlh$A2$Z$A1_EQ_1_AN_A3_EQ_0 = 1.0,
       tpllh$A3$Z$A1_EQ_0_AN_A2_EQ_0 = 1.0,
       tphhl$A3$Z$A1_EQ_0_AN_A2_EQ_0 = 1.0,
       tpllh$A3$Z$A1_EQ_1_AN_A2_EQ_1 = 1.0,
       tphhl$A3$Z$A1_EQ_1_AN_A2_EQ_1 = 1.0,
       tplhl$A3$Z$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tphlh$A3$Z$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tplhl$A3$Z$A1_EQ_1_AN_A2_EQ_0 = 1.0,
       tphlh$A3$Z$A1_EQ_1_AN_A2_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1)
       (A3 *> Z) = (tpllh$A3$Z$A1_EQ_1_AN_A2_EQ_1, tphhl$A3$Z$A1_EQ_1_AN_A2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0)
       (A3 *> Z) = (tphlh$A3$Z$A1_EQ_1_AN_A2_EQ_0, tplhl$A3$Z$A1_EQ_1_AN_A2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1)
       (A3 *> Z) = (tphlh$A3$Z$A1_EQ_0_AN_A2_EQ_1, tplhl$A3$Z$A1_EQ_0_AN_A2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0)
       (A3 *> Z) = (tpllh$A3$Z$A1_EQ_0_AN_A2_EQ_0, tphhl$A3$Z$A1_EQ_0_AN_A2_EQ_0);
     ifnone
       (A3 *> Z) = (tpllh$A3$Z,tplhl$A3$Z);

     if (A1 == 1'b1 && A3 == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_A3_EQ_1, tphhl$A2$Z$A1_EQ_1_AN_A3_EQ_1);
     if (A1 == 1'b1 && A3 == 1'b0)
       (A2 *> Z) = (tphlh$A2$Z$A1_EQ_1_AN_A3_EQ_0, tplhl$A2$Z$A1_EQ_1_AN_A3_EQ_0);
     if (A1 == 1'b0 && A3 == 1'b1)
       (A2 *> Z) = (tphlh$A2$Z$A1_EQ_0_AN_A3_EQ_1, tplhl$A2$Z$A1_EQ_0_AN_A3_EQ_1);
     if (A1 == 1'b0 && A3 == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_0_AN_A3_EQ_0, tphhl$A2$Z$A1_EQ_0_AN_A3_EQ_0);
     ifnone
       (A2 *> Z) = (tpllh$A2$Z,tplhl$A2$Z);

     if (A2 == 1'b1 && A3 == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_A3_EQ_1, tphhl$A1$Z$A2_EQ_1_AN_A3_EQ_1);
     if (A2 == 1'b1 && A3 == 1'b0)
       (A1 *> Z) = (tphlh$A1$Z$A2_EQ_1_AN_A3_EQ_0, tplhl$A1$Z$A2_EQ_1_AN_A3_EQ_0);
     if (A2 == 1'b0 && A3 == 1'b1)
       (A1 *> Z) = (tphlh$A1$Z$A2_EQ_0_AN_A3_EQ_1, tplhl$A1$Z$A2_EQ_0_AN_A3_EQ_1);
     if (A2 == 1'b0 && A3 == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_0_AN_A3_EQ_0, tphhl$A1$Z$A2_EQ_0_AN_A3_EQ_0);
     ifnone
       (A1 *> Z) = (tpllh$A1$Z,tplhl$A1$Z);*/

     // path delays
      (posedge A1 => (Z +: Z)) = (1.0, 1.0);
      (negedge A1 => (Z -: Z)) = (1.0, 1.0);
      if (A2 == 1'b1 && A3 == 1'b1) (A1 +=> Z) = (1.0, 1.0);
      if (A2 == 1'b0 && A3 == 1'b0) (A1 +=> Z) = (1.0, 1.0);
      if (A2 == 1'b0 && A3 == 1'b1) (A1 -=> Z) = (1.0, 1.0);
      if (A2 == 1'b1 && A3 == 1'b0) (A1 -=> Z) = (1.0, 1.0);


      (posedge A2 => (Z +: Z)) = (1.0, 1.0);
      (negedge A2 => (Z -: Z)) = (1.0, 1.0);
      if (A1 == 1'b1 && A3 == 1'b1) (A2 +=> Z) = (1.0, 1.0);
      if (A1 == 1'b0 && A3 == 1'b0) (A2 +=> Z) = (1.0, 1.0);
      if (A1 == 1'b0 && A3 == 1'b1) (A2 -=> Z) = (1.0, 1.0);
      if (A1 == 1'b1 && A3 == 1'b0) (A2 -=> Z) = (1.0, 1.0);


      (posedge A3 => (Z +: Z)) = (1.0, 1.0);
      (negedge A3 => (Z -: Z)) = (1.0, 1.0);
      if (A1 == 1'b0 && A2 == 1'b0) (A3 +=> Z) = (1.0, 1.0);
      if (A1 == 1'b1 && A2 == 1'b1) (A3 +=> Z) = (1.0, 1.0);
      if (A1 == 1'b0 && A2 == 1'b1) (A3 -=> Z) = (1.0, 1.0);
      if (A1 == 1'b1 && A2 == 1'b0) (A3 -=> Z) = (1.0, 1.0);



   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_XO03D2 (Z, A1, A2, A3);
input  A1 ;
input  A2 ;
input  A3 ;
output Z ;

   xor (I0_out, A1, A2);
   xor (Z, I0_out, A3);

   specify
     // delay parameters
 /*    specparam
       tpllh$A1$Z = 1.0,
       tplhl$A1$Z = 1.0,
       tphlh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tplhl$A2$Z = 1.0,
       tphlh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$A3$Z = 1.0,
       tplhl$A3$Z = 1.0,
       tphlh$A3$Z = 1.0,
       tphhl$A3$Z = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_A3_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_A3_EQ_1 = 1.0,
       tpllh$A1$Z$A2_EQ_0_AN_A3_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_0_AN_A3_EQ_0 = 1.0,
       tplhl$A1$Z$A2_EQ_0_AN_A3_EQ_1 = 1.0,
       tphlh$A1$Z$A2_EQ_0_AN_A3_EQ_1 = 1.0,
       tplhl$A1$Z$A2_EQ_1_AN_A3_EQ_0 = 1.0,
       tphlh$A1$Z$A2_EQ_1_AN_A3_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_A3_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_A3_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_0_AN_A3_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_0_AN_A3_EQ_0 = 1.0,
       tplhl$A2$Z$A1_EQ_0_AN_A3_EQ_1 = 1.0,
       tphlh$A2$Z$A1_EQ_0_AN_A3_EQ_1 = 1.0,
       tplhl$A2$Z$A1_EQ_1_AN_A3_EQ_0 = 1.0,
       tphlh$A2$Z$A1_EQ_1_AN_A3_EQ_0 = 1.0,
       tpllh$A3$Z$A1_EQ_0_AN_A2_EQ_0 = 1.0,
       tphhl$A3$Z$A1_EQ_0_AN_A2_EQ_0 = 1.0,
       tpllh$A3$Z$A1_EQ_1_AN_A2_EQ_1 = 1.0,
       tphhl$A3$Z$A1_EQ_1_AN_A2_EQ_1 = 1.0,
       tplhl$A3$Z$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tphlh$A3$Z$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tplhl$A3$Z$A1_EQ_1_AN_A2_EQ_0 = 1.0,
       tphlh$A3$Z$A1_EQ_1_AN_A2_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1)
       (A3 *> Z) = (tpllh$A3$Z$A1_EQ_1_AN_A2_EQ_1, tphhl$A3$Z$A1_EQ_1_AN_A2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0)
       (A3 *> Z) = (tphlh$A3$Z$A1_EQ_1_AN_A2_EQ_0, tplhl$A3$Z$A1_EQ_1_AN_A2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1)
       (A3 *> Z) = (tphlh$A3$Z$A1_EQ_0_AN_A2_EQ_1, tplhl$A3$Z$A1_EQ_0_AN_A2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0)
       (A3 *> Z) = (tpllh$A3$Z$A1_EQ_0_AN_A2_EQ_0, tphhl$A3$Z$A1_EQ_0_AN_A2_EQ_0);
     ifnone
       (A3 *> Z) = (tpllh$A3$Z,tplhl$A3$Z);

     if (A1 == 1'b1 && A3 == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_A3_EQ_1, tphhl$A2$Z$A1_EQ_1_AN_A3_EQ_1);
     if (A1 == 1'b1 && A3 == 1'b0)
       (A2 *> Z) = (tphlh$A2$Z$A1_EQ_1_AN_A3_EQ_0, tplhl$A2$Z$A1_EQ_1_AN_A3_EQ_0);
     if (A1 == 1'b0 && A3 == 1'b1)
       (A2 *> Z) = (tphlh$A2$Z$A1_EQ_0_AN_A3_EQ_1, tplhl$A2$Z$A1_EQ_0_AN_A3_EQ_1);
     if (A1 == 1'b0 && A3 == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_0_AN_A3_EQ_0, tphhl$A2$Z$A1_EQ_0_AN_A3_EQ_0);
     ifnone
       (A2 *> Z) = (tpllh$A2$Z,tplhl$A2$Z);

     if (A2 == 1'b1 && A3 == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_A3_EQ_1, tphhl$A1$Z$A2_EQ_1_AN_A3_EQ_1);
     if (A2 == 1'b1 && A3 == 1'b0)
       (A1 *> Z) = (tphlh$A1$Z$A2_EQ_1_AN_A3_EQ_0, tplhl$A1$Z$A2_EQ_1_AN_A3_EQ_0);
     if (A2 == 1'b0 && A3 == 1'b1)
       (A1 *> Z) = (tphlh$A1$Z$A2_EQ_0_AN_A3_EQ_1, tplhl$A1$Z$A2_EQ_0_AN_A3_EQ_1);
     if (A2 == 1'b0 && A3 == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_0_AN_A3_EQ_0, tphhl$A1$Z$A2_EQ_0_AN_A3_EQ_0);
     ifnone
       (A1 *> Z) = (tpllh$A1$Z,tplhl$A1$Z);*/

     // path delays
      (posedge A1 => (Z +: Z)) = (1.0, 1.0);
      (negedge A1 => (Z -: Z)) = (1.0, 1.0);
      if (A2 == 1'b1 && A3 == 1'b1) (A1 +=> Z) = (1.0, 1.0);
      if (A2 == 1'b0 && A3 == 1'b0) (A1 +=> Z) = (1.0, 1.0);
      if (A2 == 1'b0 && A3 == 1'b1) (A1 -=> Z) = (1.0, 1.0);
      if (A2 == 1'b1 && A3 == 1'b0) (A1 -=> Z) = (1.0, 1.0);


      (posedge A2 => (Z +: Z)) = (1.0, 1.0);
      (negedge A2 => (Z -: Z)) = (1.0, 1.0);
      if (A1 == 1'b1 && A3 == 1'b1) (A2 +=> Z) = (1.0, 1.0);
      if (A1 == 1'b0 && A3 == 1'b0) (A2 +=> Z) = (1.0, 1.0);
      if (A1 == 1'b0 && A3 == 1'b1) (A2 -=> Z) = (1.0, 1.0);
      if (A1 == 1'b1 && A3 == 1'b0) (A2 -=> Z) = (1.0, 1.0);


      (posedge A3 => (Z +: Z)) = (1.0, 1.0);
      (negedge A3 => (Z -: Z)) = (1.0, 1.0);
      if (A1 == 1'b0 && A2 == 1'b0) (A3 +=> Z) = (1.0, 1.0);
      if (A1 == 1'b1 && A2 == 1'b1) (A3 +=> Z) = (1.0, 1.0);
      if (A1 == 1'b0 && A2 == 1'b1) (A3 -=> Z) = (1.0, 1.0);
      if (A1 == 1'b1 && A2 == 1'b0) (A3 -=> Z) = (1.0, 1.0);


   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RT8_XO03D4 (Z, A1, A2, A3);
input  A1 ;
input  A2 ;
input  A3 ;
output Z ;

   xor (I0_out, A1, A2);
   xor (Z, I0_out, A3);

   specify
     // delay parameters
 /*    specparam
       tpllh$A1$Z = 1.0,
       tplhl$A1$Z = 1.0,
       tphlh$A1$Z = 1.0,
       tphhl$A1$Z = 1.0,
       tpllh$A2$Z = 1.0,
       tplhl$A2$Z = 1.0,
       tphlh$A2$Z = 1.0,
       tphhl$A2$Z = 1.0,
       tpllh$A3$Z = 1.0,
       tplhl$A3$Z = 1.0,
       tphlh$A3$Z = 1.0,
       tphhl$A3$Z = 1.0,
       tpllh$A1$Z$A2_EQ_1_AN_A3_EQ_1 = 1.0,
       tphhl$A1$Z$A2_EQ_1_AN_A3_EQ_1 = 1.0,
       tpllh$A1$Z$A2_EQ_0_AN_A3_EQ_0 = 1.0,
       tphhl$A1$Z$A2_EQ_0_AN_A3_EQ_0 = 1.0,
       tplhl$A1$Z$A2_EQ_0_AN_A3_EQ_1 = 1.0,
       tphlh$A1$Z$A2_EQ_0_AN_A3_EQ_1 = 1.0,
       tplhl$A1$Z$A2_EQ_1_AN_A3_EQ_0 = 1.0,
       tphlh$A1$Z$A2_EQ_1_AN_A3_EQ_0 = 1.0,
       tpllh$A2$Z$A1_EQ_1_AN_A3_EQ_1 = 1.0,
       tphhl$A2$Z$A1_EQ_1_AN_A3_EQ_1 = 1.0,
       tpllh$A2$Z$A1_EQ_0_AN_A3_EQ_0 = 1.0,
       tphhl$A2$Z$A1_EQ_0_AN_A3_EQ_0 = 1.0,
       tplhl$A2$Z$A1_EQ_0_AN_A3_EQ_1 = 1.0,
       tphlh$A2$Z$A1_EQ_0_AN_A3_EQ_1 = 1.0,
       tplhl$A2$Z$A1_EQ_1_AN_A3_EQ_0 = 1.0,
       tphlh$A2$Z$A1_EQ_1_AN_A3_EQ_0 = 1.0,
       tpllh$A3$Z$A1_EQ_0_AN_A2_EQ_0 = 1.0,
       tphhl$A3$Z$A1_EQ_0_AN_A2_EQ_0 = 1.0,
       tpllh$A3$Z$A1_EQ_1_AN_A2_EQ_1 = 1.0,
       tphhl$A3$Z$A1_EQ_1_AN_A2_EQ_1 = 1.0,
       tplhl$A3$Z$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tphlh$A3$Z$A1_EQ_0_AN_A2_EQ_1 = 1.0,
       tplhl$A3$Z$A1_EQ_1_AN_A2_EQ_0 = 1.0,
       tphlh$A3$Z$A1_EQ_1_AN_A2_EQ_0 = 1.0;

     // path delays
     if (A1 == 1'b1 && A2 == 1'b1)
       (A3 *> Z) = (tpllh$A3$Z$A1_EQ_1_AN_A2_EQ_1, tphhl$A3$Z$A1_EQ_1_AN_A2_EQ_1);
     if (A1 == 1'b1 && A2 == 1'b0)
       (A3 *> Z) = (tphlh$A3$Z$A1_EQ_1_AN_A2_EQ_0, tplhl$A3$Z$A1_EQ_1_AN_A2_EQ_0);
     if (A1 == 1'b0 && A2 == 1'b1)
       (A3 *> Z) = (tphlh$A3$Z$A1_EQ_0_AN_A2_EQ_1, tplhl$A3$Z$A1_EQ_0_AN_A2_EQ_1);
     if (A1 == 1'b0 && A2 == 1'b0)
       (A3 *> Z) = (tpllh$A3$Z$A1_EQ_0_AN_A2_EQ_0, tphhl$A3$Z$A1_EQ_0_AN_A2_EQ_0);
     ifnone
       (A3 *> Z) = (tpllh$A3$Z,tplhl$A3$Z);

     if (A1 == 1'b1 && A3 == 1'b1)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_1_AN_A3_EQ_1, tphhl$A2$Z$A1_EQ_1_AN_A3_EQ_1);
     if (A1 == 1'b1 && A3 == 1'b0)
       (A2 *> Z) = (tphlh$A2$Z$A1_EQ_1_AN_A3_EQ_0, tplhl$A2$Z$A1_EQ_1_AN_A3_EQ_0);
     if (A1 == 1'b0 && A3 == 1'b1)
       (A2 *> Z) = (tphlh$A2$Z$A1_EQ_0_AN_A3_EQ_1, tplhl$A2$Z$A1_EQ_0_AN_A3_EQ_1);
     if (A1 == 1'b0 && A3 == 1'b0)
       (A2 *> Z) = (tpllh$A2$Z$A1_EQ_0_AN_A3_EQ_0, tphhl$A2$Z$A1_EQ_0_AN_A3_EQ_0);
     ifnone
       (A2 *> Z) = (tpllh$A2$Z,tplhl$A2$Z);

     if (A2 == 1'b1 && A3 == 1'b1)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_1_AN_A3_EQ_1, tphhl$A1$Z$A2_EQ_1_AN_A3_EQ_1);
     if (A2 == 1'b1 && A3 == 1'b0)
       (A1 *> Z) = (tphlh$A1$Z$A2_EQ_1_AN_A3_EQ_0, tplhl$A1$Z$A2_EQ_1_AN_A3_EQ_0);
     if (A2 == 1'b0 && A3 == 1'b1)
       (A1 *> Z) = (tphlh$A1$Z$A2_EQ_0_AN_A3_EQ_1, tplhl$A1$Z$A2_EQ_0_AN_A3_EQ_1);
     if (A2 == 1'b0 && A3 == 1'b0)
       (A1 *> Z) = (tpllh$A1$Z$A2_EQ_0_AN_A3_EQ_0, tphhl$A1$Z$A2_EQ_0_AN_A3_EQ_0);
     ifnone
       (A1 *> Z) = (tpllh$A1$Z,tplhl$A1$Z);*/

  // path delays
      (posedge A1 => (Z +: Z)) = (1.0, 1.0);
      (negedge A1 => (Z -: Z)) = (1.0, 1.0);
      if (A2 == 1'b1 && A3 == 1'b1) (A1 +=> Z) = (1.0, 1.0);
      if (A2 == 1'b0 && A3 == 1'b0) (A1 +=> Z) = (1.0, 1.0);
      if (A2 == 1'b0 && A3 == 1'b1) (A1 -=> Z) = (1.0, 1.0);
      if (A2 == 1'b1 && A3 == 1'b0) (A1 -=> Z) = (1.0, 1.0);


      (posedge A2 => (Z +: Z)) = (1.0, 1.0);
      (negedge A2 => (Z -: Z)) = (1.0, 1.0);
      if (A1 == 1'b1 && A3 == 1'b1) (A2 +=> Z) = (1.0, 1.0);
      if (A1 == 1'b0 && A3 == 1'b0) (A2 +=> Z) = (1.0, 1.0);
      if (A1 == 1'b0 && A3 == 1'b1) (A2 -=> Z) = (1.0, 1.0);
      if (A1 == 1'b1 && A3 == 1'b0) (A2 -=> Z) = (1.0, 1.0);


      (posedge A3 => (Z +: Z)) = (1.0, 1.0);
      (negedge A3 => (Z -: Z)) = (1.0, 1.0);
      if (A1 == 1'b0 && A2 == 1'b0) (A3 +=> Z) = (1.0, 1.0);
      if (A1 == 1'b1 && A2 == 1'b1) (A3 +=> Z) = (1.0, 1.0);
      if (A1 == 1'b0 && A2 == 1'b1) (A3 -=> Z) = (1.0, 1.0);
      if (A1 == 1'b1 && A2 == 1'b0) (A3 -=> Z) = (1.0, 1.0);



   endspecify

endmodule
`endcelldefine

primitive udp_dff (out, in, clk, clr, set, NOTIFIER);
   output out;
   input  in, clk, clr, set, NOTIFIER;
   reg    out;

   table

// in  clk  clr   set  NOT  : Qt : Qt+1
//
   0  r   ?   0   ?   : ?  :  0  ; // clock in 0
   1  r   0   ?   ?   : ?  :  1  ; // clock in 1
   1  *   0   ?   ?   : 1  :  1  ; // reduce pessimism
   0  *   ?   0   ?   : 0  :  0  ; // reduce pessimism
   ?  f   ?   ?   ?   : ?  :  -  ; // no changes on negedge clk
   *  b   ?   ?   ?   : ?  :  -  ; // no changes when in switches
   ?  ?   ?   1   ?   : ?  :  1  ; // set output
   ?  b   0   *   ?   : 1  :  1  ; // cover all transistions on set
   1  x   0   *   ?   : 1  :  1  ; // cover all transistions on set
   ?  ?   1   0   ?   : ?  :  0  ; // reset output
   ?  b   *   0   ?   : 0  :  0  ; // cover all transistions on clr
   0  x   *   0   ?   : 0  :  0  ; // cover all transistions on clr
   ?  ?   ?   ?   *   : ?  :  x  ; // any notifier changed

   endtable
endprimitive // udp_dff

primitive udp_tlat (out, in, enable, clr, set, NOTIFIER);

   output out;
   input  in, enable, clr, set, NOTIFIER;
   reg    out;

   table

// in  enable  clr   set  NOT  : Qt : Qt+1
//
   1  1   0   ?   ?   : ?  :  1  ; //
   0  1   ?   0   ?   : ?  :  0  ; //
   1  *   0   ?   ?   : 1  :  1  ; // reduce pessimism
   0  *   ?   0   ?   : 0  :  0  ; // reduce pessimism
   *  0   ?   ?   ?   : ?  :  -  ; // no changes when in switches
   ?  ?   ?   1   ?   : ?  :  1  ; // set output
   ?  0   0   *   ?   : 1  :  1  ; // cover all transistions on set
   1  ?   0   *   ?   : 1  :  1  ; // cover all transistions on set
   ?  ?   1   0   ?   : ?  :  0  ; // reset output
   ?  0   *   0   ?   : 0  :  0  ; // cover all transistions on clr
   0  ?   *   0   ?   : 0  :  0  ; // cover all transistions on clr
   ?  ?   ?   ?   *   : ?  :  x  ; // any notifier changed

   endtable
endprimitive // udp_tlat

primitive udp_mux2 (out, in0, in1, sel);
   output out;
   input  in0, in1, sel;

   table

// in0 in1 sel :  out
//
    1  ?  0 :  1 ;
    0  ?  0 :  0 ;
    ?  1  1 :  1 ;
    ?  0  1 :  0 ;
    0  0  x :  0 ;
    1  1  x :  1 ;

   endtable
endprimitive // udp_mux2

